module background_rom(
        input wire clk,
        input wire [8:0] x,
        input wire [7:0] y,
        output reg [11:0] color_data
);

    (* rom_style = "block" *)

    //signal declaration
    reg [8:0] x_reg;
    reg [7:0] y_reg;

    always @(posedge clk) begin
        x_reg <= x;
        y_reg <= y;
    end

    always @*
        case ({x_reg, y_reg})
			// right: 9'd319, bottom: 8'd239
			{9'd0, 8'd45}: color_data = 12'h000;
			{9'd0, 8'd46}: color_data = 12'h000;
			{9'd0, 8'd47}: color_data = 12'h000;
			{9'd0, 8'd48}: color_data = 12'h000;
			{9'd0, 8'd49}: color_data = 12'h000;
			{9'd0, 8'd50}: color_data = 12'h000;
			{9'd0, 8'd51}: color_data = 12'h560;
			{9'd0, 8'd52}: color_data = 12'h9b0;
			{9'd0, 8'd53}: color_data = 12'hcd7;
			{9'd0, 8'd54}: color_data = 12'hfff;
			{9'd0, 8'd55}: color_data = 12'hdea;
			{9'd0, 8'd56}: color_data = 12'h9b0;
			{9'd0, 8'd57}: color_data = 12'h9b0;
			{9'd0, 8'd58}: color_data = 12'h9a0;
			{9'd0, 8'd59}: color_data = 12'h560;
			{9'd0, 8'd60}: color_data = 12'h020;
			{9'd0, 8'd61}: color_data = 12'h130;
			{9'd0, 8'd62}: color_data = 12'h240;
			{9'd0, 8'd63}: color_data = 12'h560;
			{9'd0, 8'd64}: color_data = 12'h760;
			{9'd0, 8'd65}: color_data = 12'h220;
			{9'd0, 8'd68}: color_data = 12'h057;
			{9'd0, 8'd69}: color_data = 12'h0cf;
			{9'd0, 8'd70}: color_data = 12'h0bf;
			{9'd0, 8'd71}: color_data = 12'h0bf;
			{9'd0, 8'd72}: color_data = 12'h0bf;
			{9'd0, 8'd73}: color_data = 12'h0bf;
			{9'd0, 8'd74}: color_data = 12'h0bf;
			{9'd0, 8'd75}: color_data = 12'h0cf;
			{9'd0, 8'd76}: color_data = 12'h0ae;
			{9'd0, 8'd77}: color_data = 12'h023;
			{9'd0, 8'd128}: color_data = 12'h057;
			{9'd0, 8'd129}: color_data = 12'h0cf;
			{9'd0, 8'd130}: color_data = 12'h0bf;
			{9'd0, 8'd131}: color_data = 12'h0bf;
			{9'd0, 8'd132}: color_data = 12'h0bf;
			{9'd0, 8'd133}: color_data = 12'h0bf;
			{9'd0, 8'd134}: color_data = 12'h0bf;
			{9'd0, 8'd135}: color_data = 12'h0bf;
			{9'd0, 8'd136}: color_data = 12'h0ae;
			{9'd0, 8'd137}: color_data = 12'h023;
			{9'd0, 8'd170}: color_data = 12'h000;
			{9'd0, 8'd171}: color_data = 12'h068;
			{9'd0, 8'd172}: color_data = 12'h0cf;
			{9'd0, 8'd173}: color_data = 12'h0bf;
			{9'd0, 8'd174}: color_data = 12'h0bf;
			{9'd0, 8'd175}: color_data = 12'h0bf;
			{9'd0, 8'd176}: color_data = 12'h0bf;
			{9'd0, 8'd177}: color_data = 12'h0bf;
			{9'd0, 8'd178}: color_data = 12'h0cf;
			{9'd0, 8'd179}: color_data = 12'h09d;
			{9'd0, 8'd180}: color_data = 12'h012;
			{9'd0, 8'd205}: color_data = 12'h330;
			{9'd0, 8'd206}: color_data = 12'h9b0;
			{9'd0, 8'd207}: color_data = 12'hbc3;
			{9'd0, 8'd208}: color_data = 12'hffe;
			{9'd0, 8'd209}: color_data = 12'hffd;
			{9'd0, 8'd210}: color_data = 12'hac2;
			{9'd0, 8'd211}: color_data = 12'h9b0;
			{9'd0, 8'd212}: color_data = 12'h9b0;
			{9'd0, 8'd213}: color_data = 12'h9b0;
			{9'd0, 8'd214}: color_data = 12'h780;
			{9'd0, 8'd215}: color_data = 12'h230;
			{9'd0, 8'd216}: color_data = 12'h030;
			{9'd0, 8'd217}: color_data = 12'h140;
			{9'd0, 8'd218}: color_data = 12'h450;
			{9'd0, 8'd219}: color_data = 12'h770;
			{9'd0, 8'd220}: color_data = 12'h440;
			{9'd0, 8'd221}: color_data = 12'h000;
			{9'd0, 8'd222}: color_data = 12'h000;
			{9'd0, 8'd223}: color_data = 12'h000;
			{9'd0, 8'd224}: color_data = 12'h000;
			{9'd0, 8'd225}: color_data = 12'h000;
			{9'd0, 8'd226}: color_data = 12'h000;
			{9'd0, 8'd227}: color_data = 12'h700;
			{9'd0, 8'd228}: color_data = 12'ha00;
			{9'd0, 8'd229}: color_data = 12'h900;
			{9'd0, 8'd230}: color_data = 12'h300;
			{9'd0, 8'd232}: color_data = 12'h000;
			{9'd0, 8'd233}: color_data = 12'h000;
			{9'd0, 8'd235}: color_data = 12'h300;
			{9'd0, 8'd236}: color_data = 12'h900;
			{9'd0, 8'd237}: color_data = 12'ha00;
			{9'd0, 8'd238}: color_data = 12'h700;
			{9'd0, 8'd239}: color_data = 12'h100;
			{9'd1, 8'd24}: color_data = 12'h000;
			{9'd1, 8'd25}: color_data = 12'h000;
			{9'd1, 8'd26}: color_data = 12'h000;
			{9'd1, 8'd27}: color_data = 12'h000;
			{9'd1, 8'd28}: color_data = 12'h000;
			{9'd1, 8'd29}: color_data = 12'h000;
			{9'd1, 8'd30}: color_data = 12'h000;
			{9'd1, 8'd31}: color_data = 12'h000;
			{9'd1, 8'd32}: color_data = 12'h000;
			{9'd1, 8'd33}: color_data = 12'h000;
			{9'd1, 8'd34}: color_data = 12'h000;
			{9'd1, 8'd35}: color_data = 12'h000;
			{9'd1, 8'd36}: color_data = 12'h000;
			{9'd1, 8'd37}: color_data = 12'h000;
			{9'd1, 8'd38}: color_data = 12'h000;
			{9'd1, 8'd39}: color_data = 12'h000;
			{9'd1, 8'd40}: color_data = 12'h000;
			{9'd1, 8'd41}: color_data = 12'h000;
			{9'd1, 8'd42}: color_data = 12'h000;
			{9'd1, 8'd43}: color_data = 12'h000;
			{9'd1, 8'd45}: color_data = 12'h111;
			{9'd1, 8'd46}: color_data = 12'h888;
			{9'd1, 8'd47}: color_data = 12'h783;
			{9'd1, 8'd48}: color_data = 12'h670;
			{9'd1, 8'd49}: color_data = 12'h670;
			{9'd1, 8'd50}: color_data = 12'h220;
			{9'd1, 8'd51}: color_data = 12'h450;
			{9'd1, 8'd52}: color_data = 12'h9b0;
			{9'd1, 8'd53}: color_data = 12'hcd7;
			{9'd1, 8'd54}: color_data = 12'hfff;
			{9'd1, 8'd55}: color_data = 12'hdea;
			{9'd1, 8'd56}: color_data = 12'h9b0;
			{9'd1, 8'd57}: color_data = 12'h9b0;
			{9'd1, 8'd58}: color_data = 12'h9a0;
			{9'd1, 8'd59}: color_data = 12'h560;
			{9'd1, 8'd60}: color_data = 12'h020;
			{9'd1, 8'd61}: color_data = 12'h130;
			{9'd1, 8'd62}: color_data = 12'h240;
			{9'd1, 8'd63}: color_data = 12'h560;
			{9'd1, 8'd64}: color_data = 12'h760;
			{9'd1, 8'd65}: color_data = 12'h220;
			{9'd1, 8'd68}: color_data = 12'h047;
			{9'd1, 8'd69}: color_data = 12'h4df;
			{9'd1, 8'd70}: color_data = 12'h7df;
			{9'd1, 8'd71}: color_data = 12'h0bf;
			{9'd1, 8'd72}: color_data = 12'h0bf;
			{9'd1, 8'd73}: color_data = 12'h0cf;
			{9'd1, 8'd74}: color_data = 12'h0ad;
			{9'd1, 8'd75}: color_data = 12'h068;
			{9'd1, 8'd76}: color_data = 12'h09c;
			{9'd1, 8'd77}: color_data = 12'h034;
			{9'd1, 8'd128}: color_data = 12'h047;
			{9'd1, 8'd129}: color_data = 12'h4df;
			{9'd1, 8'd130}: color_data = 12'h7df;
			{9'd1, 8'd131}: color_data = 12'h0bf;
			{9'd1, 8'd132}: color_data = 12'h0bf;
			{9'd1, 8'd133}: color_data = 12'h0cf;
			{9'd1, 8'd134}: color_data = 12'h0ad;
			{9'd1, 8'd135}: color_data = 12'h068;
			{9'd1, 8'd136}: color_data = 12'h09c;
			{9'd1, 8'd137}: color_data = 12'h034;
			{9'd1, 8'd170}: color_data = 12'h000;
			{9'd1, 8'd171}: color_data = 12'h068;
			{9'd1, 8'd172}: color_data = 12'h5df;
			{9'd1, 8'd173}: color_data = 12'h6df;
			{9'd1, 8'd174}: color_data = 12'h0bf;
			{9'd1, 8'd175}: color_data = 12'h0bf;
			{9'd1, 8'd176}: color_data = 12'h0cf;
			{9'd1, 8'd177}: color_data = 12'h09c;
			{9'd1, 8'd178}: color_data = 12'h068;
			{9'd1, 8'd179}: color_data = 12'h08c;
			{9'd1, 8'd180}: color_data = 12'h023;
			{9'd1, 8'd205}: color_data = 12'h330;
			{9'd1, 8'd206}: color_data = 12'h9b0;
			{9'd1, 8'd207}: color_data = 12'hbc3;
			{9'd1, 8'd208}: color_data = 12'hffe;
			{9'd1, 8'd209}: color_data = 12'hffd;
			{9'd1, 8'd210}: color_data = 12'hac2;
			{9'd1, 8'd211}: color_data = 12'h9b0;
			{9'd1, 8'd212}: color_data = 12'h9b0;
			{9'd1, 8'd213}: color_data = 12'h9b0;
			{9'd1, 8'd214}: color_data = 12'h780;
			{9'd1, 8'd215}: color_data = 12'h230;
			{9'd1, 8'd216}: color_data = 12'h030;
			{9'd1, 8'd217}: color_data = 12'h140;
			{9'd1, 8'd218}: color_data = 12'h450;
			{9'd1, 8'd219}: color_data = 12'h770;
			{9'd1, 8'd220}: color_data = 12'h440;
			{9'd1, 8'd221}: color_data = 12'h000;
			{9'd1, 8'd222}: color_data = 12'h100;
			{9'd1, 8'd223}: color_data = 12'h500;
			{9'd1, 8'd224}: color_data = 12'h600;
			{9'd1, 8'd225}: color_data = 12'h500;
			{9'd1, 8'd226}: color_data = 12'h200;
			{9'd1, 8'd227}: color_data = 12'ha20;
			{9'd1, 8'd228}: color_data = 12'hb10;
			{9'd1, 8'd229}: color_data = 12'h900;
			{9'd1, 8'd230}: color_data = 12'h300;
			{9'd1, 8'd231}: color_data = 12'h200;
			{9'd1, 8'd232}: color_data = 12'h600;
			{9'd1, 8'd233}: color_data = 12'h600;
			{9'd1, 8'd234}: color_data = 12'h200;
			{9'd1, 8'd235}: color_data = 12'h410;
			{9'd1, 8'd236}: color_data = 12'hc20;
			{9'd1, 8'd237}: color_data = 12'ha00;
			{9'd1, 8'd238}: color_data = 12'h700;
			{9'd1, 8'd239}: color_data = 12'h100;
			{9'd2, 8'd24}: color_data = 12'h120;
			{9'd2, 8'd25}: color_data = 12'h450;
			{9'd2, 8'd26}: color_data = 12'h450;
			{9'd2, 8'd27}: color_data = 12'h450;
			{9'd2, 8'd28}: color_data = 12'h450;
			{9'd2, 8'd29}: color_data = 12'h450;
			{9'd2, 8'd30}: color_data = 12'h450;
			{9'd2, 8'd31}: color_data = 12'h450;
			{9'd2, 8'd32}: color_data = 12'h450;
			{9'd2, 8'd33}: color_data = 12'h450;
			{9'd2, 8'd34}: color_data = 12'h450;
			{9'd2, 8'd35}: color_data = 12'h460;
			{9'd2, 8'd36}: color_data = 12'h460;
			{9'd2, 8'd37}: color_data = 12'h460;
			{9'd2, 8'd38}: color_data = 12'h460;
			{9'd2, 8'd39}: color_data = 12'h460;
			{9'd2, 8'd40}: color_data = 12'h460;
			{9'd2, 8'd41}: color_data = 12'h460;
			{9'd2, 8'd42}: color_data = 12'h460;
			{9'd2, 8'd43}: color_data = 12'h450;
			{9'd2, 8'd44}: color_data = 12'h450;
			{9'd2, 8'd45}: color_data = 12'h662;
			{9'd2, 8'd46}: color_data = 12'hdec;
			{9'd2, 8'd47}: color_data = 12'hbd4;
			{9'd2, 8'd48}: color_data = 12'h9c0;
			{9'd2, 8'd49}: color_data = 12'h9c0;
			{9'd2, 8'd50}: color_data = 12'h340;
			{9'd2, 8'd51}: color_data = 12'h460;
			{9'd2, 8'd52}: color_data = 12'h9b0;
			{9'd2, 8'd53}: color_data = 12'hcd7;
			{9'd2, 8'd54}: color_data = 12'hfff;
			{9'd2, 8'd55}: color_data = 12'hdea;
			{9'd2, 8'd56}: color_data = 12'h9b0;
			{9'd2, 8'd57}: color_data = 12'h9b0;
			{9'd2, 8'd58}: color_data = 12'h9a0;
			{9'd2, 8'd59}: color_data = 12'h560;
			{9'd2, 8'd60}: color_data = 12'h020;
			{9'd2, 8'd61}: color_data = 12'h130;
			{9'd2, 8'd62}: color_data = 12'h240;
			{9'd2, 8'd63}: color_data = 12'h560;
			{9'd2, 8'd64}: color_data = 12'h760;
			{9'd2, 8'd65}: color_data = 12'h220;
			{9'd2, 8'd68}: color_data = 12'h047;
			{9'd2, 8'd69}: color_data = 12'h6df;
			{9'd2, 8'd70}: color_data = 12'heff;
			{9'd2, 8'd71}: color_data = 12'h6df;
			{9'd2, 8'd72}: color_data = 12'h0bf;
			{9'd2, 8'd73}: color_data = 12'h0be;
			{9'd2, 8'd74}: color_data = 12'h056;
			{9'd2, 8'd75}: color_data = 12'h012;
			{9'd2, 8'd76}: color_data = 12'h08b;
			{9'd2, 8'd77}: color_data = 12'h034;
			{9'd2, 8'd128}: color_data = 12'h047;
			{9'd2, 8'd129}: color_data = 12'h6df;
			{9'd2, 8'd130}: color_data = 12'heff;
			{9'd2, 8'd131}: color_data = 12'h6df;
			{9'd2, 8'd132}: color_data = 12'h0bf;
			{9'd2, 8'd133}: color_data = 12'h0be;
			{9'd2, 8'd134}: color_data = 12'h056;
			{9'd2, 8'd135}: color_data = 12'h012;
			{9'd2, 8'd136}: color_data = 12'h08b;
			{9'd2, 8'd137}: color_data = 12'h034;
			{9'd2, 8'd170}: color_data = 12'h000;
			{9'd2, 8'd171}: color_data = 12'h068;
			{9'd2, 8'd172}: color_data = 12'h8ef;
			{9'd2, 8'd173}: color_data = 12'hdff;
			{9'd2, 8'd174}: color_data = 12'h4cf;
			{9'd2, 8'd175}: color_data = 12'h0bf;
			{9'd2, 8'd176}: color_data = 12'h0ae;
			{9'd2, 8'd177}: color_data = 12'h035;
			{9'd2, 8'd178}: color_data = 12'h023;
			{9'd2, 8'd179}: color_data = 12'h08c;
			{9'd2, 8'd180}: color_data = 12'h023;
			{9'd2, 8'd205}: color_data = 12'h330;
			{9'd2, 8'd206}: color_data = 12'h9b0;
			{9'd2, 8'd207}: color_data = 12'hbc3;
			{9'd2, 8'd208}: color_data = 12'hffe;
			{9'd2, 8'd209}: color_data = 12'hffd;
			{9'd2, 8'd210}: color_data = 12'hac2;
			{9'd2, 8'd211}: color_data = 12'h9b0;
			{9'd2, 8'd212}: color_data = 12'h9b0;
			{9'd2, 8'd213}: color_data = 12'h9b0;
			{9'd2, 8'd214}: color_data = 12'h780;
			{9'd2, 8'd215}: color_data = 12'h230;
			{9'd2, 8'd216}: color_data = 12'h030;
			{9'd2, 8'd217}: color_data = 12'h140;
			{9'd2, 8'd218}: color_data = 12'h450;
			{9'd2, 8'd219}: color_data = 12'h770;
			{9'd2, 8'd220}: color_data = 12'h440;
			{9'd2, 8'd221}: color_data = 12'h000;
			{9'd2, 8'd222}: color_data = 12'h200;
			{9'd2, 8'd223}: color_data = 12'h900;
			{9'd2, 8'd224}: color_data = 12'hb00;
			{9'd2, 8'd225}: color_data = 12'h800;
			{9'd2, 8'd226}: color_data = 12'h200;
			{9'd2, 8'd227}: color_data = 12'hb30;
			{9'd2, 8'd228}: color_data = 12'hc10;
			{9'd2, 8'd229}: color_data = 12'h800;
			{9'd2, 8'd230}: color_data = 12'h300;
			{9'd2, 8'd231}: color_data = 12'h400;
			{9'd2, 8'd232}: color_data = 12'ha00;
			{9'd2, 8'd233}: color_data = 12'ha00;
			{9'd2, 8'd234}: color_data = 12'h500;
			{9'd2, 8'd235}: color_data = 12'h510;
			{9'd2, 8'd236}: color_data = 12'hd30;
			{9'd2, 8'd237}: color_data = 12'ha00;
			{9'd2, 8'd238}: color_data = 12'h700;
			{9'd2, 8'd239}: color_data = 12'h100;
			{9'd3, 8'd22}: color_data = 12'h110;
			{9'd3, 8'd23}: color_data = 12'h230;
			{9'd3, 8'd24}: color_data = 12'h560;
			{9'd3, 8'd25}: color_data = 12'h9c0;
			{9'd3, 8'd26}: color_data = 12'h9b0;
			{9'd3, 8'd27}: color_data = 12'h9b0;
			{9'd3, 8'd28}: color_data = 12'h9b0;
			{9'd3, 8'd29}: color_data = 12'h9b0;
			{9'd3, 8'd30}: color_data = 12'h9b0;
			{9'd3, 8'd31}: color_data = 12'h9b0;
			{9'd3, 8'd32}: color_data = 12'h9b0;
			{9'd3, 8'd33}: color_data = 12'h9c0;
			{9'd3, 8'd34}: color_data = 12'h9c0;
			{9'd3, 8'd35}: color_data = 12'haa0;
			{9'd3, 8'd36}: color_data = 12'hc70;
			{9'd3, 8'd37}: color_data = 12'hc70;
			{9'd3, 8'd38}: color_data = 12'hc80;
			{9'd3, 8'd39}: color_data = 12'hc80;
			{9'd3, 8'd40}: color_data = 12'hc70;
			{9'd3, 8'd41}: color_data = 12'hc70;
			{9'd3, 8'd42}: color_data = 12'hb90;
			{9'd3, 8'd43}: color_data = 12'h9c0;
			{9'd3, 8'd44}: color_data = 12'h9c0;
			{9'd3, 8'd45}: color_data = 12'hac2;
			{9'd3, 8'd46}: color_data = 12'hefc;
			{9'd3, 8'd47}: color_data = 12'hde8;
			{9'd3, 8'd48}: color_data = 12'hbd4;
			{9'd3, 8'd49}: color_data = 12'hbd5;
			{9'd3, 8'd50}: color_data = 12'h462;
			{9'd3, 8'd51}: color_data = 12'h460;
			{9'd3, 8'd52}: color_data = 12'hac1;
			{9'd3, 8'd53}: color_data = 12'hdea;
			{9'd3, 8'd54}: color_data = 12'hfff;
			{9'd3, 8'd55}: color_data = 12'hdea;
			{9'd3, 8'd56}: color_data = 12'h9b0;
			{9'd3, 8'd57}: color_data = 12'h9b0;
			{9'd3, 8'd58}: color_data = 12'h9a0;
			{9'd3, 8'd59}: color_data = 12'h560;
			{9'd3, 8'd60}: color_data = 12'h020;
			{9'd3, 8'd61}: color_data = 12'h130;
			{9'd3, 8'd62}: color_data = 12'h240;
			{9'd3, 8'd63}: color_data = 12'h560;
			{9'd3, 8'd64}: color_data = 12'h760;
			{9'd3, 8'd65}: color_data = 12'h220;
			{9'd3, 8'd68}: color_data = 12'h047;
			{9'd3, 8'd69}: color_data = 12'h6df;
			{9'd3, 8'd70}: color_data = 12'hfff;
			{9'd3, 8'd71}: color_data = 12'hdff;
			{9'd3, 8'd72}: color_data = 12'h5df;
			{9'd3, 8'd73}: color_data = 12'h068;
			{9'd3, 8'd74}: color_data = 12'h000;
			{9'd3, 8'd75}: color_data = 12'h012;
			{9'd3, 8'd76}: color_data = 12'h08c;
			{9'd3, 8'd77}: color_data = 12'h034;
			{9'd3, 8'd128}: color_data = 12'h047;
			{9'd3, 8'd129}: color_data = 12'h6df;
			{9'd3, 8'd130}: color_data = 12'hfff;
			{9'd3, 8'd131}: color_data = 12'hdff;
			{9'd3, 8'd132}: color_data = 12'h5df;
			{9'd3, 8'd133}: color_data = 12'h068;
			{9'd3, 8'd134}: color_data = 12'h000;
			{9'd3, 8'd135}: color_data = 12'h012;
			{9'd3, 8'd136}: color_data = 12'h08c;
			{9'd3, 8'd137}: color_data = 12'h034;
			{9'd3, 8'd170}: color_data = 12'h000;
			{9'd3, 8'd171}: color_data = 12'h068;
			{9'd3, 8'd172}: color_data = 12'h8ef;
			{9'd3, 8'd173}: color_data = 12'hfff;
			{9'd3, 8'd174}: color_data = 12'hcff;
			{9'd3, 8'd175}: color_data = 12'h4ce;
			{9'd3, 8'd176}: color_data = 12'h057;
			{9'd3, 8'd177}: color_data = 12'h000;
			{9'd3, 8'd178}: color_data = 12'h023;
			{9'd3, 8'd179}: color_data = 12'h08c;
			{9'd3, 8'd180}: color_data = 12'h023;
			{9'd3, 8'd205}: color_data = 12'h330;
			{9'd3, 8'd206}: color_data = 12'h9b0;
			{9'd3, 8'd207}: color_data = 12'hbc3;
			{9'd3, 8'd208}: color_data = 12'hffe;
			{9'd3, 8'd209}: color_data = 12'hffd;
			{9'd3, 8'd210}: color_data = 12'hac2;
			{9'd3, 8'd211}: color_data = 12'h9b0;
			{9'd3, 8'd212}: color_data = 12'h9b0;
			{9'd3, 8'd213}: color_data = 12'h9b0;
			{9'd3, 8'd214}: color_data = 12'h780;
			{9'd3, 8'd215}: color_data = 12'h230;
			{9'd3, 8'd216}: color_data = 12'h030;
			{9'd3, 8'd217}: color_data = 12'h140;
			{9'd3, 8'd218}: color_data = 12'h450;
			{9'd3, 8'd219}: color_data = 12'h770;
			{9'd3, 8'd220}: color_data = 12'h440;
			{9'd3, 8'd221}: color_data = 12'h000;
			{9'd3, 8'd222}: color_data = 12'h200;
			{9'd3, 8'd223}: color_data = 12'h900;
			{9'd3, 8'd224}: color_data = 12'ha00;
			{9'd3, 8'd225}: color_data = 12'h700;
			{9'd3, 8'd226}: color_data = 12'h200;
			{9'd3, 8'd227}: color_data = 12'hb30;
			{9'd3, 8'd228}: color_data = 12'he20;
			{9'd3, 8'd229}: color_data = 12'ha00;
			{9'd3, 8'd230}: color_data = 12'h300;
			{9'd3, 8'd231}: color_data = 12'h400;
			{9'd3, 8'd232}: color_data = 12'ha00;
			{9'd3, 8'd233}: color_data = 12'ha00;
			{9'd3, 8'd234}: color_data = 12'h400;
			{9'd3, 8'd235}: color_data = 12'h510;
			{9'd3, 8'd236}: color_data = 12'hf40;
			{9'd3, 8'd237}: color_data = 12'hd10;
			{9'd3, 8'd238}: color_data = 12'h800;
			{9'd3, 8'd239}: color_data = 12'h100;
			{9'd4, 8'd21}: color_data = 12'h000;
			{9'd4, 8'd22}: color_data = 12'h560;
			{9'd4, 8'd23}: color_data = 12'h9b0;
			{9'd4, 8'd24}: color_data = 12'h9b0;
			{9'd4, 8'd25}: color_data = 12'h9b0;
			{9'd4, 8'd26}: color_data = 12'hac3;
			{9'd4, 8'd27}: color_data = 12'hac2;
			{9'd4, 8'd28}: color_data = 12'hac0;
			{9'd4, 8'd29}: color_data = 12'hac2;
			{9'd4, 8'd30}: color_data = 12'hac2;
			{9'd4, 8'd31}: color_data = 12'h9b0;
			{9'd4, 8'd32}: color_data = 12'h9b0;
			{9'd4, 8'd33}: color_data = 12'h9c0;
			{9'd4, 8'd34}: color_data = 12'hab0;
			{9'd4, 8'd35}: color_data = 12'he40;
			{9'd4, 8'd36}: color_data = 12'hf10;
			{9'd4, 8'd37}: color_data = 12'he20;
			{9'd4, 8'd38}: color_data = 12'hf10;
			{9'd4, 8'd39}: color_data = 12'hf10;
			{9'd4, 8'd40}: color_data = 12'he10;
			{9'd4, 8'd41}: color_data = 12'hf10;
			{9'd4, 8'd42}: color_data = 12'he20;
			{9'd4, 8'd43}: color_data = 12'ha90;
			{9'd4, 8'd44}: color_data = 12'h8b0;
			{9'd4, 8'd45}: color_data = 12'hac1;
			{9'd4, 8'd46}: color_data = 12'hefc;
			{9'd4, 8'd47}: color_data = 12'hfff;
			{9'd4, 8'd48}: color_data = 12'hfff;
			{9'd4, 8'd49}: color_data = 12'hffe;
			{9'd4, 8'd50}: color_data = 12'h565;
			{9'd4, 8'd51}: color_data = 12'h460;
			{9'd4, 8'd52}: color_data = 12'hde8;
			{9'd4, 8'd53}: color_data = 12'hfff;
			{9'd4, 8'd54}: color_data = 12'hfff;
			{9'd4, 8'd55}: color_data = 12'hdd8;
			{9'd4, 8'd56}: color_data = 12'h9b0;
			{9'd4, 8'd57}: color_data = 12'h9b0;
			{9'd4, 8'd58}: color_data = 12'h9a0;
			{9'd4, 8'd59}: color_data = 12'h560;
			{9'd4, 8'd60}: color_data = 12'h020;
			{9'd4, 8'd61}: color_data = 12'h130;
			{9'd4, 8'd62}: color_data = 12'h240;
			{9'd4, 8'd63}: color_data = 12'h560;
			{9'd4, 8'd64}: color_data = 12'h760;
			{9'd4, 8'd65}: color_data = 12'h220;
			{9'd4, 8'd68}: color_data = 12'h047;
			{9'd4, 8'd69}: color_data = 12'h6df;
			{9'd4, 8'd70}: color_data = 12'hfff;
			{9'd4, 8'd71}: color_data = 12'hfff;
			{9'd4, 8'd72}: color_data = 12'h9aa;
			{9'd4, 8'd73}: color_data = 12'h011;
			{9'd4, 8'd75}: color_data = 12'h012;
			{9'd4, 8'd76}: color_data = 12'h08c;
			{9'd4, 8'd77}: color_data = 12'h034;
			{9'd4, 8'd128}: color_data = 12'h047;
			{9'd4, 8'd129}: color_data = 12'h6df;
			{9'd4, 8'd130}: color_data = 12'hfff;
			{9'd4, 8'd131}: color_data = 12'hfff;
			{9'd4, 8'd132}: color_data = 12'h9aa;
			{9'd4, 8'd133}: color_data = 12'h111;
			{9'd4, 8'd135}: color_data = 12'h012;
			{9'd4, 8'd136}: color_data = 12'h08c;
			{9'd4, 8'd137}: color_data = 12'h034;
			{9'd4, 8'd170}: color_data = 12'h000;
			{9'd4, 8'd171}: color_data = 12'h068;
			{9'd4, 8'd172}: color_data = 12'h7ef;
			{9'd4, 8'd173}: color_data = 12'hfff;
			{9'd4, 8'd174}: color_data = 12'hfff;
			{9'd4, 8'd175}: color_data = 12'h899;
			{9'd4, 8'd176}: color_data = 12'h001;
			{9'd4, 8'd178}: color_data = 12'h024;
			{9'd4, 8'd179}: color_data = 12'h08c;
			{9'd4, 8'd180}: color_data = 12'h023;
			{9'd4, 8'd205}: color_data = 12'h330;
			{9'd4, 8'd206}: color_data = 12'h9b0;
			{9'd4, 8'd207}: color_data = 12'hbc3;
			{9'd4, 8'd208}: color_data = 12'hffe;
			{9'd4, 8'd209}: color_data = 12'hffd;
			{9'd4, 8'd210}: color_data = 12'hac2;
			{9'd4, 8'd211}: color_data = 12'h9b0;
			{9'd4, 8'd212}: color_data = 12'h9b0;
			{9'd4, 8'd213}: color_data = 12'h9b0;
			{9'd4, 8'd214}: color_data = 12'h780;
			{9'd4, 8'd215}: color_data = 12'h230;
			{9'd4, 8'd216}: color_data = 12'h030;
			{9'd4, 8'd217}: color_data = 12'h140;
			{9'd4, 8'd218}: color_data = 12'h450;
			{9'd4, 8'd219}: color_data = 12'h770;
			{9'd4, 8'd220}: color_data = 12'h440;
			{9'd4, 8'd221}: color_data = 12'h000;
			{9'd4, 8'd222}: color_data = 12'h200;
			{9'd4, 8'd223}: color_data = 12'h800;
			{9'd4, 8'd224}: color_data = 12'ha00;
			{9'd4, 8'd225}: color_data = 12'h800;
			{9'd4, 8'd226}: color_data = 12'h200;
			{9'd4, 8'd227}: color_data = 12'h920;
			{9'd4, 8'd228}: color_data = 12'hd30;
			{9'd4, 8'd229}: color_data = 12'h910;
			{9'd4, 8'd230}: color_data = 12'h200;
			{9'd4, 8'd231}: color_data = 12'h400;
			{9'd4, 8'd232}: color_data = 12'h900;
			{9'd4, 8'd233}: color_data = 12'ha00;
			{9'd4, 8'd234}: color_data = 12'h400;
			{9'd4, 8'd235}: color_data = 12'h310;
			{9'd4, 8'd236}: color_data = 12'hc30;
			{9'd4, 8'd237}: color_data = 12'hc20;
			{9'd4, 8'd238}: color_data = 12'h600;
			{9'd4, 8'd239}: color_data = 12'h000;
			{9'd5, 8'd20}: color_data = 12'h000;
			{9'd5, 8'd21}: color_data = 12'h450;
			{9'd5, 8'd22}: color_data = 12'h9b0;
			{9'd5, 8'd23}: color_data = 12'hac0;
			{9'd5, 8'd24}: color_data = 12'h9b0;
			{9'd5, 8'd25}: color_data = 12'hbc5;
			{9'd5, 8'd26}: color_data = 12'hefd;
			{9'd5, 8'd27}: color_data = 12'hde9;
			{9'd5, 8'd28}: color_data = 12'hac3;
			{9'd5, 8'd29}: color_data = 12'heeb;
			{9'd5, 8'd30}: color_data = 12'heec;
			{9'd5, 8'd31}: color_data = 12'hac2;
			{9'd5, 8'd32}: color_data = 12'h8b0;
			{9'd5, 8'd33}: color_data = 12'h9b0;
			{9'd5, 8'd34}: color_data = 12'hd40;
			{9'd5, 8'd35}: color_data = 12'hf00;
			{9'd5, 8'd36}: color_data = 12'hc50;
			{9'd5, 8'd37}: color_data = 12'h870;
			{9'd5, 8'd38}: color_data = 12'hc20;
			{9'd5, 8'd39}: color_data = 12'hd10;
			{9'd5, 8'd40}: color_data = 12'h750;
			{9'd5, 8'd41}: color_data = 12'ha30;
			{9'd5, 8'd42}: color_data = 12'hf00;
			{9'd5, 8'd43}: color_data = 12'hd20;
			{9'd5, 8'd44}: color_data = 12'h760;
			{9'd5, 8'd45}: color_data = 12'h9b1;
			{9'd5, 8'd46}: color_data = 12'hefc;
			{9'd5, 8'd47}: color_data = 12'hfff;
			{9'd5, 8'd48}: color_data = 12'hfff;
			{9'd5, 8'd49}: color_data = 12'hffe;
			{9'd5, 8'd50}: color_data = 12'h565;
			{9'd5, 8'd51}: color_data = 12'h786;
			{9'd5, 8'd52}: color_data = 12'hfff;
			{9'd5, 8'd53}: color_data = 12'hfff;
			{9'd5, 8'd54}: color_data = 12'hdea;
			{9'd5, 8'd55}: color_data = 12'hab1;
			{9'd5, 8'd56}: color_data = 12'h9b0;
			{9'd5, 8'd57}: color_data = 12'h9b0;
			{9'd5, 8'd58}: color_data = 12'h9a0;
			{9'd5, 8'd59}: color_data = 12'h560;
			{9'd5, 8'd60}: color_data = 12'h020;
			{9'd5, 8'd61}: color_data = 12'h130;
			{9'd5, 8'd62}: color_data = 12'h240;
			{9'd5, 8'd63}: color_data = 12'h560;
			{9'd5, 8'd64}: color_data = 12'h760;
			{9'd5, 8'd65}: color_data = 12'h220;
			{9'd5, 8'd68}: color_data = 12'h047;
			{9'd5, 8'd69}: color_data = 12'h6df;
			{9'd5, 8'd70}: color_data = 12'hfff;
			{9'd5, 8'd71}: color_data = 12'hcbb;
			{9'd5, 8'd72}: color_data = 12'h323;
			{9'd5, 8'd73}: color_data = 12'h002;
			{9'd5, 8'd74}: color_data = 12'h000;
			{9'd5, 8'd75}: color_data = 12'h012;
			{9'd5, 8'd76}: color_data = 12'h08c;
			{9'd5, 8'd77}: color_data = 12'h034;
			{9'd5, 8'd128}: color_data = 12'h047;
			{9'd5, 8'd129}: color_data = 12'h6df;
			{9'd5, 8'd130}: color_data = 12'hfff;
			{9'd5, 8'd131}: color_data = 12'hcbb;
			{9'd5, 8'd132}: color_data = 12'h323;
			{9'd5, 8'd133}: color_data = 12'h002;
			{9'd5, 8'd134}: color_data = 12'h000;
			{9'd5, 8'd135}: color_data = 12'h012;
			{9'd5, 8'd136}: color_data = 12'h08c;
			{9'd5, 8'd137}: color_data = 12'h034;
			{9'd5, 8'd170}: color_data = 12'h000;
			{9'd5, 8'd171}: color_data = 12'h068;
			{9'd5, 8'd172}: color_data = 12'h8ef;
			{9'd5, 8'd173}: color_data = 12'hfff;
			{9'd5, 8'd174}: color_data = 12'haaa;
			{9'd5, 8'd175}: color_data = 12'h213;
			{9'd5, 8'd176}: color_data = 12'h002;
			{9'd5, 8'd178}: color_data = 12'h023;
			{9'd5, 8'd179}: color_data = 12'h08c;
			{9'd5, 8'd180}: color_data = 12'h023;
			{9'd5, 8'd205}: color_data = 12'h330;
			{9'd5, 8'd206}: color_data = 12'h9b0;
			{9'd5, 8'd207}: color_data = 12'hbc3;
			{9'd5, 8'd208}: color_data = 12'hffe;
			{9'd5, 8'd209}: color_data = 12'hffd;
			{9'd5, 8'd210}: color_data = 12'hac2;
			{9'd5, 8'd211}: color_data = 12'h9b0;
			{9'd5, 8'd212}: color_data = 12'h9b0;
			{9'd5, 8'd213}: color_data = 12'h9b0;
			{9'd5, 8'd214}: color_data = 12'h780;
			{9'd5, 8'd215}: color_data = 12'h230;
			{9'd5, 8'd216}: color_data = 12'h030;
			{9'd5, 8'd217}: color_data = 12'h140;
			{9'd5, 8'd218}: color_data = 12'h450;
			{9'd5, 8'd219}: color_data = 12'h770;
			{9'd5, 8'd220}: color_data = 12'h440;
			{9'd5, 8'd221}: color_data = 12'h000;
			{9'd5, 8'd222}: color_data = 12'h200;
			{9'd5, 8'd223}: color_data = 12'h900;
			{9'd5, 8'd224}: color_data = 12'ha00;
			{9'd5, 8'd225}: color_data = 12'h800;
			{9'd5, 8'd226}: color_data = 12'h100;
			{9'd5, 8'd227}: color_data = 12'h100;
			{9'd5, 8'd228}: color_data = 12'h310;
			{9'd5, 8'd229}: color_data = 12'h200;
			{9'd5, 8'd230}: color_data = 12'h000;
			{9'd5, 8'd231}: color_data = 12'h500;
			{9'd5, 8'd232}: color_data = 12'ha00;
			{9'd5, 8'd233}: color_data = 12'ha00;
			{9'd5, 8'd234}: color_data = 12'h500;
			{9'd5, 8'd235}: color_data = 12'h000;
			{9'd5, 8'd236}: color_data = 12'h200;
			{9'd5, 8'd237}: color_data = 12'h300;
			{9'd5, 8'd238}: color_data = 12'h100;
			{9'd5, 8'd239}: color_data = 12'h000;
			{9'd6, 8'd19}: color_data = 12'h000;
			{9'd6, 8'd20}: color_data = 12'h340;
			{9'd6, 8'd21}: color_data = 12'h8a0;
			{9'd6, 8'd22}: color_data = 12'h9b0;
			{9'd6, 8'd23}: color_data = 12'hbc4;
			{9'd6, 8'd24}: color_data = 12'hdea;
			{9'd6, 8'd25}: color_data = 12'hefc;
			{9'd6, 8'd26}: color_data = 12'hfff;
			{9'd6, 8'd27}: color_data = 12'heeb;
			{9'd6, 8'd28}: color_data = 12'hac3;
			{9'd6, 8'd29}: color_data = 12'hffd;
			{9'd6, 8'd30}: color_data = 12'hffe;
			{9'd6, 8'd31}: color_data = 12'hac3;
			{9'd6, 8'd32}: color_data = 12'h9b0;
			{9'd6, 8'd33}: color_data = 12'hc50;
			{9'd6, 8'd34}: color_data = 12'hf00;
			{9'd6, 8'd35}: color_data = 12'hd40;
			{9'd6, 8'd36}: color_data = 12'h890;
			{9'd6, 8'd37}: color_data = 12'h6a0;
			{9'd6, 8'd38}: color_data = 12'hb50;
			{9'd6, 8'd39}: color_data = 12'hd30;
			{9'd6, 8'd40}: color_data = 12'h690;
			{9'd6, 8'd41}: color_data = 12'h680;
			{9'd6, 8'd42}: color_data = 12'hc50;
			{9'd6, 8'd43}: color_data = 12'hf00;
			{9'd6, 8'd44}: color_data = 12'hc10;
			{9'd6, 8'd45}: color_data = 12'h882;
			{9'd6, 8'd46}: color_data = 12'hdec;
			{9'd6, 8'd47}: color_data = 12'hde8;
			{9'd6, 8'd48}: color_data = 12'hbd4;
			{9'd6, 8'd49}: color_data = 12'hbc5;
			{9'd6, 8'd50}: color_data = 12'h351;
			{9'd6, 8'd51}: color_data = 12'h898;
			{9'd6, 8'd52}: color_data = 12'hfff;
			{9'd6, 8'd53}: color_data = 12'heeb;
			{9'd6, 8'd54}: color_data = 12'hac2;
			{9'd6, 8'd55}: color_data = 12'h9b0;
			{9'd6, 8'd56}: color_data = 12'h9b0;
			{9'd6, 8'd57}: color_data = 12'h9b0;
			{9'd6, 8'd58}: color_data = 12'h9a0;
			{9'd6, 8'd59}: color_data = 12'h560;
			{9'd6, 8'd60}: color_data = 12'h020;
			{9'd6, 8'd61}: color_data = 12'h130;
			{9'd6, 8'd62}: color_data = 12'h240;
			{9'd6, 8'd63}: color_data = 12'h560;
			{9'd6, 8'd64}: color_data = 12'h760;
			{9'd6, 8'd65}: color_data = 12'h220;
			{9'd6, 8'd68}: color_data = 12'h047;
			{9'd6, 8'd69}: color_data = 12'h6ef;
			{9'd6, 8'd70}: color_data = 12'hdcc;
			{9'd6, 8'd71}: color_data = 12'h434;
			{9'd6, 8'd72}: color_data = 12'h003;
			{9'd6, 8'd73}: color_data = 12'h005;
			{9'd6, 8'd74}: color_data = 12'h002;
			{9'd6, 8'd75}: color_data = 12'h012;
			{9'd6, 8'd76}: color_data = 12'h08c;
			{9'd6, 8'd77}: color_data = 12'h034;
			{9'd6, 8'd128}: color_data = 12'h047;
			{9'd6, 8'd129}: color_data = 12'h6ef;
			{9'd6, 8'd130}: color_data = 12'hddc;
			{9'd6, 8'd131}: color_data = 12'h434;
			{9'd6, 8'd132}: color_data = 12'h003;
			{9'd6, 8'd133}: color_data = 12'h005;
			{9'd6, 8'd134}: color_data = 12'h002;
			{9'd6, 8'd135}: color_data = 12'h012;
			{9'd6, 8'd136}: color_data = 12'h08c;
			{9'd6, 8'd137}: color_data = 12'h034;
			{9'd6, 8'd170}: color_data = 12'h000;
			{9'd6, 8'd171}: color_data = 12'h068;
			{9'd6, 8'd172}: color_data = 12'h8ff;
			{9'd6, 8'd173}: color_data = 12'hcbb;
			{9'd6, 8'd174}: color_data = 12'h323;
			{9'd6, 8'd175}: color_data = 12'h003;
			{9'd6, 8'd176}: color_data = 12'h005;
			{9'd6, 8'd177}: color_data = 12'h002;
			{9'd6, 8'd178}: color_data = 12'h023;
			{9'd6, 8'd179}: color_data = 12'h09c;
			{9'd6, 8'd180}: color_data = 12'h023;
			{9'd6, 8'd205}: color_data = 12'h330;
			{9'd6, 8'd206}: color_data = 12'h9b0;
			{9'd6, 8'd207}: color_data = 12'hbc3;
			{9'd6, 8'd208}: color_data = 12'hffe;
			{9'd6, 8'd209}: color_data = 12'hffd;
			{9'd6, 8'd210}: color_data = 12'hac2;
			{9'd6, 8'd211}: color_data = 12'h9b0;
			{9'd6, 8'd212}: color_data = 12'h9b0;
			{9'd6, 8'd213}: color_data = 12'h9b0;
			{9'd6, 8'd214}: color_data = 12'h780;
			{9'd6, 8'd215}: color_data = 12'h230;
			{9'd6, 8'd216}: color_data = 12'h030;
			{9'd6, 8'd217}: color_data = 12'h140;
			{9'd6, 8'd218}: color_data = 12'h450;
			{9'd6, 8'd219}: color_data = 12'h770;
			{9'd6, 8'd220}: color_data = 12'h440;
			{9'd6, 8'd221}: color_data = 12'h000;
			{9'd6, 8'd222}: color_data = 12'h300;
			{9'd6, 8'd223}: color_data = 12'hc20;
			{9'd6, 8'd224}: color_data = 12'ha00;
			{9'd6, 8'd225}: color_data = 12'h800;
			{9'd6, 8'd226}: color_data = 12'h100;
			{9'd6, 8'd227}: color_data = 12'h300;
			{9'd6, 8'd228}: color_data = 12'h500;
			{9'd6, 8'd229}: color_data = 12'h500;
			{9'd6, 8'd230}: color_data = 12'h100;
			{9'd6, 8'd231}: color_data = 12'h710;
			{9'd6, 8'd232}: color_data = 12'hc10;
			{9'd6, 8'd233}: color_data = 12'h900;
			{9'd6, 8'd234}: color_data = 12'h500;
			{9'd6, 8'd235}: color_data = 12'h100;
			{9'd6, 8'd236}: color_data = 12'h500;
			{9'd6, 8'd237}: color_data = 12'h500;
			{9'd6, 8'd238}: color_data = 12'h400;
			{9'd6, 8'd239}: color_data = 12'h000;
			{9'd7, 8'd19}: color_data = 12'h330;
			{9'd7, 8'd20}: color_data = 12'h8a0;
			{9'd7, 8'd21}: color_data = 12'h9c0;
			{9'd7, 8'd22}: color_data = 12'hac3;
			{9'd7, 8'd23}: color_data = 12'heec;
			{9'd7, 8'd24}: color_data = 12'hfff;
			{9'd7, 8'd25}: color_data = 12'hfff;
			{9'd7, 8'd26}: color_data = 12'hffe;
			{9'd7, 8'd27}: color_data = 12'hbd5;
			{9'd7, 8'd28}: color_data = 12'hab1;
			{9'd7, 8'd29}: color_data = 12'hcd7;
			{9'd7, 8'd30}: color_data = 12'hcd7;
			{9'd7, 8'd31}: color_data = 12'h9c1;
			{9'd7, 8'd32}: color_data = 12'h9a0;
			{9'd7, 8'd33}: color_data = 12'he20;
			{9'd7, 8'd34}: color_data = 12'he30;
			{9'd7, 8'd35}: color_data = 12'h980;
			{9'd7, 8'd36}: color_data = 12'h790;
			{9'd7, 8'd37}: color_data = 12'h8b0;
			{9'd7, 8'd38}: color_data = 12'hc60;
			{9'd7, 8'd39}: color_data = 12'hd40;
			{9'd7, 8'd40}: color_data = 12'h8a0;
			{9'd7, 8'd41}: color_data = 12'h680;
			{9'd7, 8'd42}: color_data = 12'h9a0;
			{9'd7, 8'd43}: color_data = 12'hd40;
			{9'd7, 8'd44}: color_data = 12'he00;
			{9'd7, 8'd45}: color_data = 12'ha82;
			{9'd7, 8'd46}: color_data = 12'hdec;
			{9'd7, 8'd47}: color_data = 12'hbc4;
			{9'd7, 8'd48}: color_data = 12'h8b0;
			{9'd7, 8'd49}: color_data = 12'h8b0;
			{9'd7, 8'd50}: color_data = 12'h250;
			{9'd7, 8'd51}: color_data = 12'h564;
			{9'd7, 8'd52}: color_data = 12'hcd8;
			{9'd7, 8'd53}: color_data = 12'hbc4;
			{9'd7, 8'd54}: color_data = 12'h8b0;
			{9'd7, 8'd55}: color_data = 12'h9b0;
			{9'd7, 8'd56}: color_data = 12'h9b0;
			{9'd7, 8'd57}: color_data = 12'h9b0;
			{9'd7, 8'd58}: color_data = 12'h9a0;
			{9'd7, 8'd59}: color_data = 12'h560;
			{9'd7, 8'd60}: color_data = 12'h020;
			{9'd7, 8'd61}: color_data = 12'h130;
			{9'd7, 8'd62}: color_data = 12'h240;
			{9'd7, 8'd63}: color_data = 12'h560;
			{9'd7, 8'd64}: color_data = 12'h760;
			{9'd7, 8'd65}: color_data = 12'h220;
			{9'd7, 8'd68}: color_data = 12'h057;
			{9'd7, 8'd69}: color_data = 12'h3bd;
			{9'd7, 8'd70}: color_data = 12'h555;
			{9'd7, 8'd71}: color_data = 12'h002;
			{9'd7, 8'd72}: color_data = 12'h005;
			{9'd7, 8'd73}: color_data = 12'h005;
			{9'd7, 8'd74}: color_data = 12'h004;
			{9'd7, 8'd75}: color_data = 12'h025;
			{9'd7, 8'd76}: color_data = 12'h09c;
			{9'd7, 8'd77}: color_data = 12'h034;
			{9'd7, 8'd128}: color_data = 12'h057;
			{9'd7, 8'd129}: color_data = 12'h3bd;
			{9'd7, 8'd130}: color_data = 12'h555;
			{9'd7, 8'd131}: color_data = 12'h002;
			{9'd7, 8'd132}: color_data = 12'h005;
			{9'd7, 8'd133}: color_data = 12'h005;
			{9'd7, 8'd134}: color_data = 12'h004;
			{9'd7, 8'd135}: color_data = 12'h025;
			{9'd7, 8'd136}: color_data = 12'h09c;
			{9'd7, 8'd137}: color_data = 12'h034;
			{9'd7, 8'd170}: color_data = 12'h000;
			{9'd7, 8'd171}: color_data = 12'h079;
			{9'd7, 8'd172}: color_data = 12'h4bd;
			{9'd7, 8'd173}: color_data = 12'h444;
			{9'd7, 8'd174}: color_data = 12'h002;
			{9'd7, 8'd175}: color_data = 12'h005;
			{9'd7, 8'd176}: color_data = 12'h005;
			{9'd7, 8'd177}: color_data = 12'h004;
			{9'd7, 8'd178}: color_data = 12'h036;
			{9'd7, 8'd179}: color_data = 12'h09c;
			{9'd7, 8'd180}: color_data = 12'h023;
			{9'd7, 8'd205}: color_data = 12'h330;
			{9'd7, 8'd206}: color_data = 12'h9b0;
			{9'd7, 8'd207}: color_data = 12'hbc3;
			{9'd7, 8'd208}: color_data = 12'hffe;
			{9'd7, 8'd209}: color_data = 12'hffd;
			{9'd7, 8'd210}: color_data = 12'hac2;
			{9'd7, 8'd211}: color_data = 12'h9b0;
			{9'd7, 8'd212}: color_data = 12'h9b0;
			{9'd7, 8'd213}: color_data = 12'h9b0;
			{9'd7, 8'd214}: color_data = 12'h780;
			{9'd7, 8'd215}: color_data = 12'h230;
			{9'd7, 8'd216}: color_data = 12'h030;
			{9'd7, 8'd217}: color_data = 12'h140;
			{9'd7, 8'd218}: color_data = 12'h450;
			{9'd7, 8'd219}: color_data = 12'h770;
			{9'd7, 8'd220}: color_data = 12'h440;
			{9'd7, 8'd221}: color_data = 12'h000;
			{9'd7, 8'd222}: color_data = 12'h410;
			{9'd7, 8'd223}: color_data = 12'hd30;
			{9'd7, 8'd224}: color_data = 12'hb00;
			{9'd7, 8'd225}: color_data = 12'h700;
			{9'd7, 8'd226}: color_data = 12'h200;
			{9'd7, 8'd227}: color_data = 12'h700;
			{9'd7, 8'd228}: color_data = 12'hb00;
			{9'd7, 8'd229}: color_data = 12'h900;
			{9'd7, 8'd230}: color_data = 12'h300;
			{9'd7, 8'd231}: color_data = 12'h820;
			{9'd7, 8'd232}: color_data = 12'hd20;
			{9'd7, 8'd233}: color_data = 12'h900;
			{9'd7, 8'd234}: color_data = 12'h500;
			{9'd7, 8'd235}: color_data = 12'h300;
			{9'd7, 8'd236}: color_data = 12'h900;
			{9'd7, 8'd237}: color_data = 12'hb00;
			{9'd7, 8'd238}: color_data = 12'h800;
			{9'd7, 8'd239}: color_data = 12'h100;
			{9'd8, 8'd18}: color_data = 12'h220;
			{9'd8, 8'd19}: color_data = 12'h790;
			{9'd8, 8'd20}: color_data = 12'h9c0;
			{9'd8, 8'd21}: color_data = 12'hac2;
			{9'd8, 8'd22}: color_data = 12'hdea;
			{9'd8, 8'd23}: color_data = 12'hfff;
			{9'd8, 8'd24}: color_data = 12'hffe;
			{9'd8, 8'd25}: color_data = 12'heeb;
			{9'd8, 8'd26}: color_data = 12'hcd7;
			{9'd8, 8'd27}: color_data = 12'h9b0;
			{9'd8, 8'd28}: color_data = 12'h9b0;
			{9'd8, 8'd29}: color_data = 12'h9b0;
			{9'd8, 8'd30}: color_data = 12'h9b0;
			{9'd8, 8'd31}: color_data = 12'h9b0;
			{9'd8, 8'd32}: color_data = 12'h9a0;
			{9'd8, 8'd33}: color_data = 12'he30;
			{9'd8, 8'd34}: color_data = 12'hb70;
			{9'd8, 8'd35}: color_data = 12'h690;
			{9'd8, 8'd36}: color_data = 12'h7a0;
			{9'd8, 8'd37}: color_data = 12'haa0;
			{9'd8, 8'd38}: color_data = 12'he30;
			{9'd8, 8'd39}: color_data = 12'he20;
			{9'd8, 8'd40}: color_data = 12'h970;
			{9'd8, 8'd41}: color_data = 12'h680;
			{9'd8, 8'd42}: color_data = 12'h8d0;
			{9'd8, 8'd43}: color_data = 12'haa0;
			{9'd8, 8'd44}: color_data = 12'he20;
			{9'd8, 8'd45}: color_data = 12'hba2;
			{9'd8, 8'd46}: color_data = 12'hefc;
			{9'd8, 8'd47}: color_data = 12'hbc4;
			{9'd8, 8'd48}: color_data = 12'h9b0;
			{9'd8, 8'd49}: color_data = 12'h9b0;
			{9'd8, 8'd50}: color_data = 12'h350;
			{9'd8, 8'd51}: color_data = 12'h230;
			{9'd8, 8'd52}: color_data = 12'h880;
			{9'd8, 8'd53}: color_data = 12'h9b0;
			{9'd8, 8'd54}: color_data = 12'h9b0;
			{9'd8, 8'd55}: color_data = 12'h9b0;
			{9'd8, 8'd56}: color_data = 12'h9b0;
			{9'd8, 8'd57}: color_data = 12'h9b0;
			{9'd8, 8'd58}: color_data = 12'h9b0;
			{9'd8, 8'd59}: color_data = 12'h660;
			{9'd8, 8'd60}: color_data = 12'h020;
			{9'd8, 8'd61}: color_data = 12'h130;
			{9'd8, 8'd62}: color_data = 12'h240;
			{9'd8, 8'd63}: color_data = 12'h560;
			{9'd8, 8'd64}: color_data = 12'h760;
			{9'd8, 8'd65}: color_data = 12'h220;
			{9'd8, 8'd68}: color_data = 12'h036;
			{9'd8, 8'd69}: color_data = 12'h047;
			{9'd8, 8'd70}: color_data = 12'h001;
			{9'd8, 8'd71}: color_data = 12'h004;
			{9'd8, 8'd72}: color_data = 12'h004;
			{9'd8, 8'd73}: color_data = 12'h004;
			{9'd8, 8'd74}: color_data = 12'h004;
			{9'd8, 8'd75}: color_data = 12'h015;
			{9'd8, 8'd76}: color_data = 12'h059;
			{9'd8, 8'd77}: color_data = 12'h023;
			{9'd8, 8'd128}: color_data = 12'h035;
			{9'd8, 8'd129}: color_data = 12'h047;
			{9'd8, 8'd130}: color_data = 12'h001;
			{9'd8, 8'd131}: color_data = 12'h004;
			{9'd8, 8'd132}: color_data = 12'h004;
			{9'd8, 8'd133}: color_data = 12'h004;
			{9'd8, 8'd134}: color_data = 12'h004;
			{9'd8, 8'd135}: color_data = 12'h015;
			{9'd8, 8'd136}: color_data = 12'h059;
			{9'd8, 8'd137}: color_data = 12'h023;
			{9'd8, 8'd170}: color_data = 12'h000;
			{9'd8, 8'd171}: color_data = 12'h047;
			{9'd8, 8'd172}: color_data = 12'h036;
			{9'd8, 8'd173}: color_data = 12'h001;
			{9'd8, 8'd174}: color_data = 12'h004;
			{9'd8, 8'd175}: color_data = 12'h004;
			{9'd8, 8'd176}: color_data = 12'h004;
			{9'd8, 8'd177}: color_data = 12'h004;
			{9'd8, 8'd178}: color_data = 12'h016;
			{9'd8, 8'd179}: color_data = 12'h059;
			{9'd8, 8'd180}: color_data = 12'h012;
			{9'd8, 8'd205}: color_data = 12'h330;
			{9'd8, 8'd206}: color_data = 12'h9b0;
			{9'd8, 8'd207}: color_data = 12'hbc3;
			{9'd8, 8'd208}: color_data = 12'hffe;
			{9'd8, 8'd209}: color_data = 12'hffd;
			{9'd8, 8'd210}: color_data = 12'hac2;
			{9'd8, 8'd211}: color_data = 12'h9b0;
			{9'd8, 8'd212}: color_data = 12'h9b0;
			{9'd8, 8'd213}: color_data = 12'h9b0;
			{9'd8, 8'd214}: color_data = 12'h780;
			{9'd8, 8'd215}: color_data = 12'h230;
			{9'd8, 8'd216}: color_data = 12'h030;
			{9'd8, 8'd217}: color_data = 12'h140;
			{9'd8, 8'd218}: color_data = 12'h450;
			{9'd8, 8'd219}: color_data = 12'h770;
			{9'd8, 8'd220}: color_data = 12'h440;
			{9'd8, 8'd221}: color_data = 12'h000;
			{9'd8, 8'd222}: color_data = 12'h410;
			{9'd8, 8'd223}: color_data = 12'he40;
			{9'd8, 8'd224}: color_data = 12'hd20;
			{9'd8, 8'd225}: color_data = 12'h800;
			{9'd8, 8'd226}: color_data = 12'h200;
			{9'd8, 8'd227}: color_data = 12'h600;
			{9'd8, 8'd228}: color_data = 12'ha00;
			{9'd8, 8'd229}: color_data = 12'h900;
			{9'd8, 8'd230}: color_data = 12'h300;
			{9'd8, 8'd231}: color_data = 12'h820;
			{9'd8, 8'd232}: color_data = 12'hf30;
			{9'd8, 8'd233}: color_data = 12'hc00;
			{9'd8, 8'd234}: color_data = 12'h500;
			{9'd8, 8'd235}: color_data = 12'h200;
			{9'd8, 8'd236}: color_data = 12'h900;
			{9'd8, 8'd237}: color_data = 12'ha00;
			{9'd8, 8'd238}: color_data = 12'h700;
			{9'd8, 8'd239}: color_data = 12'h100;
			{9'd9, 8'd17}: color_data = 12'h000;
			{9'd9, 8'd18}: color_data = 12'h670;
			{9'd9, 8'd19}: color_data = 12'hac0;
			{9'd9, 8'd20}: color_data = 12'hac1;
			{9'd9, 8'd21}: color_data = 12'hde9;
			{9'd9, 8'd22}: color_data = 12'hfff;
			{9'd9, 8'd23}: color_data = 12'hfff;
			{9'd9, 8'd24}: color_data = 12'hcd8;
			{9'd9, 8'd25}: color_data = 12'h9b1;
			{9'd9, 8'd26}: color_data = 12'h9b0;
			{9'd9, 8'd27}: color_data = 12'h9b0;
			{9'd9, 8'd28}: color_data = 12'h9b0;
			{9'd9, 8'd29}: color_data = 12'h9b0;
			{9'd9, 8'd30}: color_data = 12'h9b0;
			{9'd9, 8'd31}: color_data = 12'h9c0;
			{9'd9, 8'd32}: color_data = 12'h9b0;
			{9'd9, 8'd33}: color_data = 12'he30;
			{9'd9, 8'd34}: color_data = 12'hc50;
			{9'd9, 8'd35}: color_data = 12'h870;
			{9'd9, 8'd36}: color_data = 12'h970;
			{9'd9, 8'd37}: color_data = 12'hd50;
			{9'd9, 8'd38}: color_data = 12'hf11;
			{9'd9, 8'd39}: color_data = 12'hf22;
			{9'd9, 8'd40}: color_data = 12'hd10;
			{9'd9, 8'd41}: color_data = 12'h960;
			{9'd9, 8'd42}: color_data = 12'haa0;
			{9'd9, 8'd43}: color_data = 12'hc70;
			{9'd9, 8'd44}: color_data = 12'he20;
			{9'd9, 8'd45}: color_data = 12'hb92;
			{9'd9, 8'd46}: color_data = 12'hdfc;
			{9'd9, 8'd47}: color_data = 12'hbc4;
			{9'd9, 8'd48}: color_data = 12'h9b0;
			{9'd9, 8'd49}: color_data = 12'h9b0;
			{9'd9, 8'd50}: color_data = 12'h350;
			{9'd9, 8'd51}: color_data = 12'h230;
			{9'd9, 8'd52}: color_data = 12'h890;
			{9'd9, 8'd53}: color_data = 12'h9c0;
			{9'd9, 8'd54}: color_data = 12'h9b0;
			{9'd9, 8'd55}: color_data = 12'h9b0;
			{9'd9, 8'd56}: color_data = 12'h9b0;
			{9'd9, 8'd57}: color_data = 12'h9b0;
			{9'd9, 8'd58}: color_data = 12'h8a0;
			{9'd9, 8'd59}: color_data = 12'h450;
			{9'd9, 8'd60}: color_data = 12'h120;
			{9'd9, 8'd61}: color_data = 12'h130;
			{9'd9, 8'd62}: color_data = 12'h240;
			{9'd9, 8'd63}: color_data = 12'h560;
			{9'd9, 8'd64}: color_data = 12'h770;
			{9'd9, 8'd65}: color_data = 12'h220;
			{9'd9, 8'd68}: color_data = 12'h013;
			{9'd9, 8'd69}: color_data = 12'h027;
			{9'd9, 8'd70}: color_data = 12'h016;
			{9'd9, 8'd71}: color_data = 12'h027;
			{9'd9, 8'd72}: color_data = 12'h027;
			{9'd9, 8'd73}: color_data = 12'h026;
			{9'd9, 8'd74}: color_data = 12'h027;
			{9'd9, 8'd75}: color_data = 12'h028;
			{9'd9, 8'd76}: color_data = 12'h027;
			{9'd9, 8'd77}: color_data = 12'h001;
			{9'd9, 8'd128}: color_data = 12'h013;
			{9'd9, 8'd129}: color_data = 12'h027;
			{9'd9, 8'd130}: color_data = 12'h016;
			{9'd9, 8'd131}: color_data = 12'h027;
			{9'd9, 8'd132}: color_data = 12'h027;
			{9'd9, 8'd133}: color_data = 12'h027;
			{9'd9, 8'd134}: color_data = 12'h027;
			{9'd9, 8'd135}: color_data = 12'h028;
			{9'd9, 8'd136}: color_data = 12'h027;
			{9'd9, 8'd137}: color_data = 12'h001;
			{9'd9, 8'd170}: color_data = 12'h000;
			{9'd9, 8'd171}: color_data = 12'h014;
			{9'd9, 8'd172}: color_data = 12'h027;
			{9'd9, 8'd173}: color_data = 12'h016;
			{9'd9, 8'd174}: color_data = 12'h027;
			{9'd9, 8'd175}: color_data = 12'h027;
			{9'd9, 8'd176}: color_data = 12'h026;
			{9'd9, 8'd177}: color_data = 12'h027;
			{9'd9, 8'd178}: color_data = 12'h028;
			{9'd9, 8'd179}: color_data = 12'h026;
			{9'd9, 8'd180}: color_data = 12'h001;
			{9'd9, 8'd205}: color_data = 12'h330;
			{9'd9, 8'd206}: color_data = 12'h9b0;
			{9'd9, 8'd207}: color_data = 12'hbc3;
			{9'd9, 8'd208}: color_data = 12'hffe;
			{9'd9, 8'd209}: color_data = 12'hffd;
			{9'd9, 8'd210}: color_data = 12'hac2;
			{9'd9, 8'd211}: color_data = 12'h9b0;
			{9'd9, 8'd212}: color_data = 12'h9b0;
			{9'd9, 8'd213}: color_data = 12'h9b0;
			{9'd9, 8'd214}: color_data = 12'h780;
			{9'd9, 8'd215}: color_data = 12'h230;
			{9'd9, 8'd216}: color_data = 12'h030;
			{9'd9, 8'd217}: color_data = 12'h140;
			{9'd9, 8'd218}: color_data = 12'h450;
			{9'd9, 8'd219}: color_data = 12'h770;
			{9'd9, 8'd220}: color_data = 12'h440;
			{9'd9, 8'd221}: color_data = 12'h000;
			{9'd9, 8'd222}: color_data = 12'h200;
			{9'd9, 8'd223}: color_data = 12'hc30;
			{9'd9, 8'd224}: color_data = 12'hc30;
			{9'd9, 8'd225}: color_data = 12'h700;
			{9'd9, 8'd226}: color_data = 12'h100;
			{9'd9, 8'd227}: color_data = 12'h600;
			{9'd9, 8'd228}: color_data = 12'ha00;
			{9'd9, 8'd229}: color_data = 12'h900;
			{9'd9, 8'd230}: color_data = 12'h300;
			{9'd9, 8'd231}: color_data = 12'h620;
			{9'd9, 8'd232}: color_data = 12'hd40;
			{9'd9, 8'd233}: color_data = 12'ha20;
			{9'd9, 8'd234}: color_data = 12'h300;
			{9'd9, 8'd235}: color_data = 12'h200;
			{9'd9, 8'd236}: color_data = 12'h900;
			{9'd9, 8'd237}: color_data = 12'ha00;
			{9'd9, 8'd238}: color_data = 12'h700;
			{9'd9, 8'd239}: color_data = 12'h100;
			{9'd10, 8'd17}: color_data = 12'h110;
			{9'd10, 8'd18}: color_data = 12'h780;
			{9'd10, 8'd19}: color_data = 12'hac0;
			{9'd10, 8'd20}: color_data = 12'hcd7;
			{9'd10, 8'd21}: color_data = 12'hfff;
			{9'd10, 8'd22}: color_data = 12'hfff;
			{9'd10, 8'd23}: color_data = 12'hde9;
			{9'd10, 8'd24}: color_data = 12'h9b1;
			{9'd10, 8'd25}: color_data = 12'h8b0;
			{9'd10, 8'd26}: color_data = 12'h9b0;
			{9'd10, 8'd27}: color_data = 12'h9b0;
			{9'd10, 8'd28}: color_data = 12'h9b0;
			{9'd10, 8'd29}: color_data = 12'h9b0;
			{9'd10, 8'd30}: color_data = 12'h9b0;
			{9'd10, 8'd31}: color_data = 12'h9b0;
			{9'd10, 8'd32}: color_data = 12'h9b0;
			{9'd10, 8'd33}: color_data = 12'he30;
			{9'd10, 8'd34}: color_data = 12'hf00;
			{9'd10, 8'd35}: color_data = 12'he10;
			{9'd10, 8'd36}: color_data = 12'he10;
			{9'd10, 8'd37}: color_data = 12'hf00;
			{9'd10, 8'd38}: color_data = 12'hf66;
			{9'd10, 8'd39}: color_data = 12'hf88;
			{9'd10, 8'd40}: color_data = 12'hf00;
			{9'd10, 8'd41}: color_data = 12'he10;
			{9'd10, 8'd42}: color_data = 12'he20;
			{9'd10, 8'd43}: color_data = 12'hf10;
			{9'd10, 8'd44}: color_data = 12'he00;
			{9'd10, 8'd45}: color_data = 12'h972;
			{9'd10, 8'd46}: color_data = 12'hdec;
			{9'd10, 8'd47}: color_data = 12'hbd4;
			{9'd10, 8'd48}: color_data = 12'h9b0;
			{9'd10, 8'd49}: color_data = 12'h9b0;
			{9'd10, 8'd50}: color_data = 12'h350;
			{9'd10, 8'd51}: color_data = 12'h330;
			{9'd10, 8'd52}: color_data = 12'h890;
			{9'd10, 8'd53}: color_data = 12'h9b0;
			{9'd10, 8'd54}: color_data = 12'h9b0;
			{9'd10, 8'd55}: color_data = 12'h9b0;
			{9'd10, 8'd56}: color_data = 12'h9b0;
			{9'd10, 8'd57}: color_data = 12'h9a0;
			{9'd10, 8'd58}: color_data = 12'h560;
			{9'd10, 8'd59}: color_data = 12'h130;
			{9'd10, 8'd60}: color_data = 12'h130;
			{9'd10, 8'd61}: color_data = 12'h140;
			{9'd10, 8'd62}: color_data = 12'h240;
			{9'd10, 8'd63}: color_data = 12'h560;
			{9'd10, 8'd64}: color_data = 12'h660;
			{9'd10, 8'd65}: color_data = 12'h220;
			{9'd10, 8'd68}: color_data = 12'h035;
			{9'd10, 8'd69}: color_data = 12'h09e;
			{9'd10, 8'd70}: color_data = 12'h09e;
			{9'd10, 8'd71}: color_data = 12'h09e;
			{9'd10, 8'd72}: color_data = 12'h09e;
			{9'd10, 8'd73}: color_data = 12'h09e;
			{9'd10, 8'd74}: color_data = 12'h09e;
			{9'd10, 8'd75}: color_data = 12'h09e;
			{9'd10, 8'd76}: color_data = 12'h08c;
			{9'd10, 8'd77}: color_data = 12'h023;
			{9'd10, 8'd128}: color_data = 12'h035;
			{9'd10, 8'd129}: color_data = 12'h09e;
			{9'd10, 8'd130}: color_data = 12'h09e;
			{9'd10, 8'd131}: color_data = 12'h09e;
			{9'd10, 8'd132}: color_data = 12'h09e;
			{9'd10, 8'd133}: color_data = 12'h09e;
			{9'd10, 8'd134}: color_data = 12'h09e;
			{9'd10, 8'd135}: color_data = 12'h09e;
			{9'd10, 8'd136}: color_data = 12'h08c;
			{9'd10, 8'd137}: color_data = 12'h023;
			{9'd10, 8'd170}: color_data = 12'h000;
			{9'd10, 8'd171}: color_data = 12'h057;
			{9'd10, 8'd172}: color_data = 12'h0ae;
			{9'd10, 8'd173}: color_data = 12'h09e;
			{9'd10, 8'd174}: color_data = 12'h09e;
			{9'd10, 8'd175}: color_data = 12'h09e;
			{9'd10, 8'd176}: color_data = 12'h09e;
			{9'd10, 8'd177}: color_data = 12'h09e;
			{9'd10, 8'd178}: color_data = 12'h09e;
			{9'd10, 8'd179}: color_data = 12'h07b;
			{9'd10, 8'd180}: color_data = 12'h012;
			{9'd10, 8'd205}: color_data = 12'h330;
			{9'd10, 8'd206}: color_data = 12'h9b0;
			{9'd10, 8'd207}: color_data = 12'hbd3;
			{9'd10, 8'd208}: color_data = 12'hffe;
			{9'd10, 8'd209}: color_data = 12'hffd;
			{9'd10, 8'd210}: color_data = 12'hac2;
			{9'd10, 8'd211}: color_data = 12'h9b0;
			{9'd10, 8'd212}: color_data = 12'h9b0;
			{9'd10, 8'd213}: color_data = 12'h9b0;
			{9'd10, 8'd214}: color_data = 12'h780;
			{9'd10, 8'd215}: color_data = 12'h230;
			{9'd10, 8'd216}: color_data = 12'h030;
			{9'd10, 8'd217}: color_data = 12'h140;
			{9'd10, 8'd218}: color_data = 12'h450;
			{9'd10, 8'd219}: color_data = 12'h770;
			{9'd10, 8'd220}: color_data = 12'h440;
			{9'd10, 8'd221}: color_data = 12'h000;
			{9'd10, 8'd222}: color_data = 12'h000;
			{9'd10, 8'd223}: color_data = 12'h200;
			{9'd10, 8'd224}: color_data = 12'h300;
			{9'd10, 8'd225}: color_data = 12'h100;
			{9'd10, 8'd226}: color_data = 12'h000;
			{9'd10, 8'd227}: color_data = 12'h700;
			{9'd10, 8'd228}: color_data = 12'ha00;
			{9'd10, 8'd229}: color_data = 12'h900;
			{9'd10, 8'd230}: color_data = 12'h300;
			{9'd10, 8'd231}: color_data = 12'h100;
			{9'd10, 8'd232}: color_data = 12'h310;
			{9'd10, 8'd233}: color_data = 12'h200;
			{9'd10, 8'd234}: color_data = 12'h000;
			{9'd10, 8'd235}: color_data = 12'h300;
			{9'd10, 8'd236}: color_data = 12'h900;
			{9'd10, 8'd237}: color_data = 12'ha00;
			{9'd10, 8'd238}: color_data = 12'h700;
			{9'd10, 8'd239}: color_data = 12'h100;
			{9'd11, 8'd16}: color_data = 12'h000;
			{9'd11, 8'd17}: color_data = 12'h560;
			{9'd11, 8'd18}: color_data = 12'h8a0;
			{9'd11, 8'd19}: color_data = 12'h9b0;
			{9'd11, 8'd20}: color_data = 12'hdea;
			{9'd11, 8'd21}: color_data = 12'hfff;
			{9'd11, 8'd22}: color_data = 12'hdeb;
			{9'd11, 8'd23}: color_data = 12'hac2;
			{9'd11, 8'd24}: color_data = 12'h9b0;
			{9'd11, 8'd25}: color_data = 12'h9b0;
			{9'd11, 8'd26}: color_data = 12'h9b0;
			{9'd11, 8'd27}: color_data = 12'h9b0;
			{9'd11, 8'd28}: color_data = 12'h9b0;
			{9'd11, 8'd29}: color_data = 12'h9b0;
			{9'd11, 8'd30}: color_data = 12'h780;
			{9'd11, 8'd31}: color_data = 12'h780;
			{9'd11, 8'd32}: color_data = 12'h870;
			{9'd11, 8'd33}: color_data = 12'hd20;
			{9'd11, 8'd34}: color_data = 12'hc20;
			{9'd11, 8'd35}: color_data = 12'h940;
			{9'd11, 8'd36}: color_data = 12'ha40;
			{9'd11, 8'd37}: color_data = 12'hc10;
			{9'd11, 8'd38}: color_data = 12'hf33;
			{9'd11, 8'd39}: color_data = 12'hf34;
			{9'd11, 8'd40}: color_data = 12'he10;
			{9'd11, 8'd41}: color_data = 12'ha30;
			{9'd11, 8'd42}: color_data = 12'h940;
			{9'd11, 8'd43}: color_data = 12'hb20;
			{9'd11, 8'd44}: color_data = 12'hd00;
			{9'd11, 8'd45}: color_data = 12'h962;
			{9'd11, 8'd46}: color_data = 12'hdec;
			{9'd11, 8'd47}: color_data = 12'hbd4;
			{9'd11, 8'd48}: color_data = 12'h9b0;
			{9'd11, 8'd49}: color_data = 12'h9b0;
			{9'd11, 8'd50}: color_data = 12'h350;
			{9'd11, 8'd51}: color_data = 12'h330;
			{9'd11, 8'd52}: color_data = 12'h770;
			{9'd11, 8'd53}: color_data = 12'h780;
			{9'd11, 8'd54}: color_data = 12'h780;
			{9'd11, 8'd55}: color_data = 12'h780;
			{9'd11, 8'd56}: color_data = 12'h880;
			{9'd11, 8'd57}: color_data = 12'h670;
			{9'd11, 8'd58}: color_data = 12'h130;
			{9'd11, 8'd59}: color_data = 12'h030;
			{9'd11, 8'd60}: color_data = 12'h140;
			{9'd11, 8'd61}: color_data = 12'h240;
			{9'd11, 8'd62}: color_data = 12'h450;
			{9'd11, 8'd63}: color_data = 12'h660;
			{9'd11, 8'd64}: color_data = 12'h330;
			{9'd11, 8'd65}: color_data = 12'h000;
			{9'd11, 8'd68}: color_data = 12'h057;
			{9'd11, 8'd69}: color_data = 12'h4ef;
			{9'd11, 8'd70}: color_data = 12'h7ef;
			{9'd11, 8'd71}: color_data = 12'h0cf;
			{9'd11, 8'd72}: color_data = 12'h0cf;
			{9'd11, 8'd73}: color_data = 12'h0df;
			{9'd11, 8'd74}: color_data = 12'h0bd;
			{9'd11, 8'd75}: color_data = 12'h068;
			{9'd11, 8'd76}: color_data = 12'h09c;
			{9'd11, 8'd77}: color_data = 12'h034;
			{9'd11, 8'd128}: color_data = 12'h057;
			{9'd11, 8'd129}: color_data = 12'h4ef;
			{9'd11, 8'd130}: color_data = 12'h7ef;
			{9'd11, 8'd131}: color_data = 12'h0cf;
			{9'd11, 8'd132}: color_data = 12'h0cf;
			{9'd11, 8'd133}: color_data = 12'h0df;
			{9'd11, 8'd134}: color_data = 12'h0bd;
			{9'd11, 8'd135}: color_data = 12'h068;
			{9'd11, 8'd136}: color_data = 12'h09c;
			{9'd11, 8'd137}: color_data = 12'h034;
			{9'd11, 8'd170}: color_data = 12'h000;
			{9'd11, 8'd171}: color_data = 12'h069;
			{9'd11, 8'd172}: color_data = 12'h6ef;
			{9'd11, 8'd173}: color_data = 12'h6ef;
			{9'd11, 8'd174}: color_data = 12'h0cf;
			{9'd11, 8'd175}: color_data = 12'h0cf;
			{9'd11, 8'd176}: color_data = 12'h0df;
			{9'd11, 8'd177}: color_data = 12'h0ac;
			{9'd11, 8'd178}: color_data = 12'h079;
			{9'd11, 8'd179}: color_data = 12'h09c;
			{9'd11, 8'd180}: color_data = 12'h023;
			{9'd11, 8'd205}: color_data = 12'h330;
			{9'd11, 8'd206}: color_data = 12'h9b0;
			{9'd11, 8'd207}: color_data = 12'hbd3;
			{9'd11, 8'd208}: color_data = 12'hffe;
			{9'd11, 8'd209}: color_data = 12'hffd;
			{9'd11, 8'd210}: color_data = 12'hac2;
			{9'd11, 8'd211}: color_data = 12'h9b0;
			{9'd11, 8'd212}: color_data = 12'h9b0;
			{9'd11, 8'd213}: color_data = 12'h9b0;
			{9'd11, 8'd214}: color_data = 12'h780;
			{9'd11, 8'd215}: color_data = 12'h230;
			{9'd11, 8'd216}: color_data = 12'h030;
			{9'd11, 8'd217}: color_data = 12'h140;
			{9'd11, 8'd218}: color_data = 12'h450;
			{9'd11, 8'd219}: color_data = 12'h770;
			{9'd11, 8'd220}: color_data = 12'h440;
			{9'd11, 8'd221}: color_data = 12'h000;
			{9'd11, 8'd222}: color_data = 12'h100;
			{9'd11, 8'd223}: color_data = 12'h400;
			{9'd11, 8'd224}: color_data = 12'h500;
			{9'd11, 8'd225}: color_data = 12'h400;
			{9'd11, 8'd226}: color_data = 12'h200;
			{9'd11, 8'd227}: color_data = 12'ha20;
			{9'd11, 8'd228}: color_data = 12'hb10;
			{9'd11, 8'd229}: color_data = 12'h900;
			{9'd11, 8'd230}: color_data = 12'h300;
			{9'd11, 8'd231}: color_data = 12'h200;
			{9'd11, 8'd232}: color_data = 12'h500;
			{9'd11, 8'd233}: color_data = 12'h500;
			{9'd11, 8'd234}: color_data = 12'h200;
			{9'd11, 8'd235}: color_data = 12'h410;
			{9'd11, 8'd236}: color_data = 12'hc20;
			{9'd11, 8'd237}: color_data = 12'ha00;
			{9'd11, 8'd238}: color_data = 12'h700;
			{9'd11, 8'd239}: color_data = 12'h100;
			{9'd12, 8'd16}: color_data = 12'h010;
			{9'd12, 8'd17}: color_data = 12'h790;
			{9'd12, 8'd18}: color_data = 12'hac0;
			{9'd12, 8'd19}: color_data = 12'hbc5;
			{9'd12, 8'd20}: color_data = 12'hefd;
			{9'd12, 8'd21}: color_data = 12'hfff;
			{9'd12, 8'd22}: color_data = 12'hcd8;
			{9'd12, 8'd23}: color_data = 12'h8b0;
			{9'd12, 8'd24}: color_data = 12'h9b0;
			{9'd12, 8'd25}: color_data = 12'h9b0;
			{9'd12, 8'd26}: color_data = 12'h9b0;
			{9'd12, 8'd27}: color_data = 12'h9b0;
			{9'd12, 8'd28}: color_data = 12'h9b0;
			{9'd12, 8'd29}: color_data = 12'h780;
			{9'd12, 8'd30}: color_data = 12'h340;
			{9'd12, 8'd31}: color_data = 12'h230;
			{9'd12, 8'd32}: color_data = 12'h330;
			{9'd12, 8'd33}: color_data = 12'hc10;
			{9'd12, 8'd34}: color_data = 12'h730;
			{9'd12, 8'd35}: color_data = 12'h150;
			{9'd12, 8'd36}: color_data = 12'h240;
			{9'd12, 8'd37}: color_data = 12'h420;
			{9'd12, 8'd38}: color_data = 12'hc00;
			{9'd12, 8'd39}: color_data = 12'hd00;
			{9'd12, 8'd40}: color_data = 12'h620;
			{9'd12, 8'd41}: color_data = 12'h240;
			{9'd12, 8'd42}: color_data = 12'h150;
			{9'd12, 8'd43}: color_data = 12'h430;
			{9'd12, 8'd44}: color_data = 12'hc00;
			{9'd12, 8'd45}: color_data = 12'h742;
			{9'd12, 8'd46}: color_data = 12'hcdc;
			{9'd12, 8'd47}: color_data = 12'hbb4;
			{9'd12, 8'd48}: color_data = 12'h890;
			{9'd12, 8'd49}: color_data = 12'h890;
			{9'd12, 8'd50}: color_data = 12'h340;
			{9'd12, 8'd51}: color_data = 12'h120;
			{9'd12, 8'd52}: color_data = 12'h340;
			{9'd12, 8'd53}: color_data = 12'h230;
			{9'd12, 8'd54}: color_data = 12'h230;
			{9'd12, 8'd55}: color_data = 12'h230;
			{9'd12, 8'd56}: color_data = 12'h330;
			{9'd12, 8'd57}: color_data = 12'h230;
			{9'd12, 8'd58}: color_data = 12'h130;
			{9'd12, 8'd59}: color_data = 12'h140;
			{9'd12, 8'd60}: color_data = 12'h240;
			{9'd12, 8'd61}: color_data = 12'h350;
			{9'd12, 8'd62}: color_data = 12'h660;
			{9'd12, 8'd63}: color_data = 12'h760;
			{9'd12, 8'd64}: color_data = 12'h220;
			{9'd12, 8'd68}: color_data = 12'h047;
			{9'd12, 8'd69}: color_data = 12'h6df;
			{9'd12, 8'd70}: color_data = 12'heff;
			{9'd12, 8'd71}: color_data = 12'h6df;
			{9'd12, 8'd72}: color_data = 12'h0bf;
			{9'd12, 8'd73}: color_data = 12'h0bf;
			{9'd12, 8'd74}: color_data = 12'h056;
			{9'd12, 8'd75}: color_data = 12'h012;
			{9'd12, 8'd76}: color_data = 12'h08b;
			{9'd12, 8'd77}: color_data = 12'h034;
			{9'd12, 8'd128}: color_data = 12'h047;
			{9'd12, 8'd129}: color_data = 12'h6df;
			{9'd12, 8'd130}: color_data = 12'heff;
			{9'd12, 8'd131}: color_data = 12'h6df;
			{9'd12, 8'd132}: color_data = 12'h0bf;
			{9'd12, 8'd133}: color_data = 12'h0bf;
			{9'd12, 8'd134}: color_data = 12'h056;
			{9'd12, 8'd135}: color_data = 12'h012;
			{9'd12, 8'd136}: color_data = 12'h08b;
			{9'd12, 8'd137}: color_data = 12'h034;
			{9'd12, 8'd170}: color_data = 12'h000;
			{9'd12, 8'd171}: color_data = 12'h068;
			{9'd12, 8'd172}: color_data = 12'h8ef;
			{9'd12, 8'd173}: color_data = 12'hdff;
			{9'd12, 8'd174}: color_data = 12'h4cf;
			{9'd12, 8'd175}: color_data = 12'h0bf;
			{9'd12, 8'd176}: color_data = 12'h0ae;
			{9'd12, 8'd177}: color_data = 12'h035;
			{9'd12, 8'd178}: color_data = 12'h023;
			{9'd12, 8'd179}: color_data = 12'h08c;
			{9'd12, 8'd180}: color_data = 12'h023;
			{9'd12, 8'd205}: color_data = 12'h230;
			{9'd12, 8'd206}: color_data = 12'h780;
			{9'd12, 8'd207}: color_data = 12'hab3;
			{9'd12, 8'd208}: color_data = 12'hfff;
			{9'd12, 8'd209}: color_data = 12'hffd;
			{9'd12, 8'd210}: color_data = 12'h9a2;
			{9'd12, 8'd211}: color_data = 12'h780;
			{9'd12, 8'd212}: color_data = 12'h890;
			{9'd12, 8'd213}: color_data = 12'h890;
			{9'd12, 8'd214}: color_data = 12'h770;
			{9'd12, 8'd215}: color_data = 12'h230;
			{9'd12, 8'd216}: color_data = 12'h030;
			{9'd12, 8'd217}: color_data = 12'h240;
			{9'd12, 8'd218}: color_data = 12'h450;
			{9'd12, 8'd219}: color_data = 12'h770;
			{9'd12, 8'd220}: color_data = 12'h440;
			{9'd12, 8'd221}: color_data = 12'h000;
			{9'd12, 8'd222}: color_data = 12'h200;
			{9'd12, 8'd223}: color_data = 12'h900;
			{9'd12, 8'd224}: color_data = 12'hb00;
			{9'd12, 8'd225}: color_data = 12'h800;
			{9'd12, 8'd226}: color_data = 12'h200;
			{9'd12, 8'd227}: color_data = 12'hb30;
			{9'd12, 8'd228}: color_data = 12'hc10;
			{9'd12, 8'd229}: color_data = 12'h800;
			{9'd12, 8'd230}: color_data = 12'h300;
			{9'd12, 8'd231}: color_data = 12'h400;
			{9'd12, 8'd232}: color_data = 12'ha00;
			{9'd12, 8'd233}: color_data = 12'ha00;
			{9'd12, 8'd234}: color_data = 12'h500;
			{9'd12, 8'd235}: color_data = 12'h510;
			{9'd12, 8'd236}: color_data = 12'hd30;
			{9'd12, 8'd237}: color_data = 12'ha00;
			{9'd12, 8'd238}: color_data = 12'h700;
			{9'd12, 8'd239}: color_data = 12'h100;
			{9'd13, 8'd16}: color_data = 12'h010;
			{9'd13, 8'd17}: color_data = 12'h780;
			{9'd13, 8'd18}: color_data = 12'hac0;
			{9'd13, 8'd19}: color_data = 12'hdea;
			{9'd13, 8'd20}: color_data = 12'hfff;
			{9'd13, 8'd21}: color_data = 12'hefd;
			{9'd13, 8'd22}: color_data = 12'hbc5;
			{9'd13, 8'd23}: color_data = 12'h9b0;
			{9'd13, 8'd24}: color_data = 12'h9b0;
			{9'd13, 8'd25}: color_data = 12'h9b0;
			{9'd13, 8'd26}: color_data = 12'h9b0;
			{9'd13, 8'd27}: color_data = 12'h9b0;
			{9'd13, 8'd28}: color_data = 12'h890;
			{9'd13, 8'd29}: color_data = 12'h440;
			{9'd13, 8'd30}: color_data = 12'h020;
			{9'd13, 8'd31}: color_data = 12'h020;
			{9'd13, 8'd32}: color_data = 12'h120;
			{9'd13, 8'd33}: color_data = 12'hc00;
			{9'd13, 8'd34}: color_data = 12'h900;
			{9'd13, 8'd35}: color_data = 12'h120;
			{9'd13, 8'd36}: color_data = 12'h030;
			{9'd13, 8'd37}: color_data = 12'h030;
			{9'd13, 8'd38}: color_data = 12'h810;
			{9'd13, 8'd39}: color_data = 12'ha10;
			{9'd13, 8'd40}: color_data = 12'h020;
			{9'd13, 8'd41}: color_data = 12'h030;
			{9'd13, 8'd42}: color_data = 12'h020;
			{9'd13, 8'd43}: color_data = 12'h710;
			{9'd13, 8'd44}: color_data = 12'hc00;
			{9'd13, 8'd45}: color_data = 12'h431;
			{9'd13, 8'd46}: color_data = 12'hac8;
			{9'd13, 8'd47}: color_data = 12'h773;
			{9'd13, 8'd48}: color_data = 12'h340;
			{9'd13, 8'd49}: color_data = 12'h440;
			{9'd13, 8'd50}: color_data = 12'h130;
			{9'd13, 8'd51}: color_data = 12'h020;
			{9'd13, 8'd52}: color_data = 12'h020;
			{9'd13, 8'd53}: color_data = 12'h020;
			{9'd13, 8'd54}: color_data = 12'h020;
			{9'd13, 8'd55}: color_data = 12'h020;
			{9'd13, 8'd56}: color_data = 12'h020;
			{9'd13, 8'd57}: color_data = 12'h030;
			{9'd13, 8'd58}: color_data = 12'h140;
			{9'd13, 8'd59}: color_data = 12'h140;
			{9'd13, 8'd60}: color_data = 12'h350;
			{9'd13, 8'd61}: color_data = 12'h660;
			{9'd13, 8'd62}: color_data = 12'h770;
			{9'd13, 8'd63}: color_data = 12'h550;
			{9'd13, 8'd64}: color_data = 12'h110;
			{9'd13, 8'd68}: color_data = 12'h047;
			{9'd13, 8'd69}: color_data = 12'h6df;
			{9'd13, 8'd70}: color_data = 12'hfff;
			{9'd13, 8'd71}: color_data = 12'hdff;
			{9'd13, 8'd72}: color_data = 12'h5df;
			{9'd13, 8'd73}: color_data = 12'h068;
			{9'd13, 8'd74}: color_data = 12'h000;
			{9'd13, 8'd75}: color_data = 12'h012;
			{9'd13, 8'd76}: color_data = 12'h08c;
			{9'd13, 8'd77}: color_data = 12'h034;
			{9'd13, 8'd128}: color_data = 12'h047;
			{9'd13, 8'd129}: color_data = 12'h6df;
			{9'd13, 8'd130}: color_data = 12'hfff;
			{9'd13, 8'd131}: color_data = 12'hdff;
			{9'd13, 8'd132}: color_data = 12'h5df;
			{9'd13, 8'd133}: color_data = 12'h069;
			{9'd13, 8'd134}: color_data = 12'h000;
			{9'd13, 8'd135}: color_data = 12'h012;
			{9'd13, 8'd136}: color_data = 12'h08c;
			{9'd13, 8'd137}: color_data = 12'h034;
			{9'd13, 8'd170}: color_data = 12'h000;
			{9'd13, 8'd171}: color_data = 12'h068;
			{9'd13, 8'd172}: color_data = 12'h8ef;
			{9'd13, 8'd173}: color_data = 12'hfff;
			{9'd13, 8'd174}: color_data = 12'hcff;
			{9'd13, 8'd175}: color_data = 12'h4ce;
			{9'd13, 8'd176}: color_data = 12'h057;
			{9'd13, 8'd177}: color_data = 12'h000;
			{9'd13, 8'd178}: color_data = 12'h023;
			{9'd13, 8'd179}: color_data = 12'h08c;
			{9'd13, 8'd180}: color_data = 12'h023;
			{9'd13, 8'd205}: color_data = 12'h110;
			{9'd13, 8'd206}: color_data = 12'h330;
			{9'd13, 8'd207}: color_data = 12'h452;
			{9'd13, 8'd208}: color_data = 12'h9a9;
			{9'd13, 8'd209}: color_data = 12'h9a9;
			{9'd13, 8'd210}: color_data = 12'h451;
			{9'd13, 8'd211}: color_data = 12'h330;
			{9'd13, 8'd212}: color_data = 12'h340;
			{9'd13, 8'd213}: color_data = 12'h340;
			{9'd13, 8'd214}: color_data = 12'h340;
			{9'd13, 8'd215}: color_data = 12'h120;
			{9'd13, 8'd216}: color_data = 12'h020;
			{9'd13, 8'd217}: color_data = 12'h130;
			{9'd13, 8'd218}: color_data = 12'h240;
			{9'd13, 8'd219}: color_data = 12'h450;
			{9'd13, 8'd220}: color_data = 12'h230;
			{9'd13, 8'd221}: color_data = 12'h000;
			{9'd13, 8'd222}: color_data = 12'h200;
			{9'd13, 8'd223}: color_data = 12'h900;
			{9'd13, 8'd224}: color_data = 12'ha00;
			{9'd13, 8'd225}: color_data = 12'h700;
			{9'd13, 8'd226}: color_data = 12'h200;
			{9'd13, 8'd227}: color_data = 12'hb30;
			{9'd13, 8'd228}: color_data = 12'he20;
			{9'd13, 8'd229}: color_data = 12'ha00;
			{9'd13, 8'd230}: color_data = 12'h300;
			{9'd13, 8'd231}: color_data = 12'h400;
			{9'd13, 8'd232}: color_data = 12'ha00;
			{9'd13, 8'd233}: color_data = 12'ha00;
			{9'd13, 8'd234}: color_data = 12'h400;
			{9'd13, 8'd235}: color_data = 12'h510;
			{9'd13, 8'd236}: color_data = 12'hf40;
			{9'd13, 8'd237}: color_data = 12'hd10;
			{9'd13, 8'd238}: color_data = 12'h800;
			{9'd13, 8'd239}: color_data = 12'h100;
			{9'd14, 8'd16}: color_data = 12'h010;
			{9'd14, 8'd17}: color_data = 12'h780;
			{9'd14, 8'd18}: color_data = 12'hac0;
			{9'd14, 8'd19}: color_data = 12'hdea;
			{9'd14, 8'd20}: color_data = 12'hfff;
			{9'd14, 8'd21}: color_data = 12'hcd7;
			{9'd14, 8'd22}: color_data = 12'h9b0;
			{9'd14, 8'd23}: color_data = 12'h9b0;
			{9'd14, 8'd24}: color_data = 12'h9b0;
			{9'd14, 8'd25}: color_data = 12'h9b0;
			{9'd14, 8'd26}: color_data = 12'h9b0;
			{9'd14, 8'd27}: color_data = 12'h8a0;
			{9'd14, 8'd28}: color_data = 12'h450;
			{9'd14, 8'd29}: color_data = 12'h020;
			{9'd14, 8'd30}: color_data = 12'h130;
			{9'd14, 8'd31}: color_data = 12'h140;
			{9'd14, 8'd32}: color_data = 12'h140;
			{9'd14, 8'd33}: color_data = 12'ha10;
			{9'd14, 8'd34}: color_data = 12'hf00;
			{9'd14, 8'd35}: color_data = 12'h820;
			{9'd14, 8'd36}: color_data = 12'h140;
			{9'd14, 8'd37}: color_data = 12'h040;
			{9'd14, 8'd38}: color_data = 12'h820;
			{9'd14, 8'd39}: color_data = 12'ha10;
			{9'd14, 8'd40}: color_data = 12'h040;
			{9'd14, 8'd41}: color_data = 12'h040;
			{9'd14, 8'd42}: color_data = 12'h620;
			{9'd14, 8'd43}: color_data = 12'he00;
			{9'd14, 8'd44}: color_data = 12'hb00;
			{9'd14, 8'd45}: color_data = 12'h440;
			{9'd14, 8'd46}: color_data = 12'h7a0;
			{9'd14, 8'd47}: color_data = 12'h350;
			{9'd14, 8'd48}: color_data = 12'h010;
			{9'd14, 8'd49}: color_data = 12'h020;
			{9'd14, 8'd50}: color_data = 12'h020;
			{9'd14, 8'd51}: color_data = 12'h030;
			{9'd14, 8'd52}: color_data = 12'h140;
			{9'd14, 8'd53}: color_data = 12'h140;
			{9'd14, 8'd54}: color_data = 12'h140;
			{9'd14, 8'd55}: color_data = 12'h140;
			{9'd14, 8'd56}: color_data = 12'h140;
			{9'd14, 8'd57}: color_data = 12'h140;
			{9'd14, 8'd58}: color_data = 12'h240;
			{9'd14, 8'd59}: color_data = 12'h350;
			{9'd14, 8'd60}: color_data = 12'h560;
			{9'd14, 8'd61}: color_data = 12'h770;
			{9'd14, 8'd62}: color_data = 12'h550;
			{9'd14, 8'd63}: color_data = 12'h110;
			{9'd14, 8'd68}: color_data = 12'h047;
			{9'd14, 8'd69}: color_data = 12'h6df;
			{9'd14, 8'd70}: color_data = 12'hfff;
			{9'd14, 8'd71}: color_data = 12'hfff;
			{9'd14, 8'd72}: color_data = 12'h9aa;
			{9'd14, 8'd73}: color_data = 12'h011;
			{9'd14, 8'd75}: color_data = 12'h012;
			{9'd14, 8'd76}: color_data = 12'h08c;
			{9'd14, 8'd77}: color_data = 12'h034;
			{9'd14, 8'd128}: color_data = 12'h047;
			{9'd14, 8'd129}: color_data = 12'h6df;
			{9'd14, 8'd130}: color_data = 12'hfff;
			{9'd14, 8'd131}: color_data = 12'hfff;
			{9'd14, 8'd132}: color_data = 12'h9aa;
			{9'd14, 8'd133}: color_data = 12'h111;
			{9'd14, 8'd135}: color_data = 12'h012;
			{9'd14, 8'd136}: color_data = 12'h08c;
			{9'd14, 8'd137}: color_data = 12'h034;
			{9'd14, 8'd170}: color_data = 12'h000;
			{9'd14, 8'd171}: color_data = 12'h068;
			{9'd14, 8'd172}: color_data = 12'h7ef;
			{9'd14, 8'd173}: color_data = 12'hfff;
			{9'd14, 8'd174}: color_data = 12'hfff;
			{9'd14, 8'd175}: color_data = 12'h899;
			{9'd14, 8'd176}: color_data = 12'h001;
			{9'd14, 8'd178}: color_data = 12'h024;
			{9'd14, 8'd179}: color_data = 12'h08c;
			{9'd14, 8'd180}: color_data = 12'h023;
			{9'd14, 8'd204}: color_data = 12'h000;
			{9'd14, 8'd205}: color_data = 12'h120;
			{9'd14, 8'd206}: color_data = 12'h230;
			{9'd14, 8'd207}: color_data = 12'h242;
			{9'd14, 8'd208}: color_data = 12'h343;
			{9'd14, 8'd209}: color_data = 12'h241;
			{9'd14, 8'd210}: color_data = 12'h130;
			{9'd14, 8'd211}: color_data = 12'h130;
			{9'd14, 8'd212}: color_data = 12'h130;
			{9'd14, 8'd213}: color_data = 12'h130;
			{9'd14, 8'd214}: color_data = 12'h130;
			{9'd14, 8'd215}: color_data = 12'h130;
			{9'd14, 8'd216}: color_data = 12'h020;
			{9'd14, 8'd217}: color_data = 12'h020;
			{9'd14, 8'd218}: color_data = 12'h020;
			{9'd14, 8'd219}: color_data = 12'h020;
			{9'd14, 8'd220}: color_data = 12'h120;
			{9'd14, 8'd221}: color_data = 12'h000;
			{9'd14, 8'd222}: color_data = 12'h200;
			{9'd14, 8'd223}: color_data = 12'h800;
			{9'd14, 8'd224}: color_data = 12'ha00;
			{9'd14, 8'd225}: color_data = 12'h800;
			{9'd14, 8'd226}: color_data = 12'h200;
			{9'd14, 8'd227}: color_data = 12'h930;
			{9'd14, 8'd228}: color_data = 12'hd30;
			{9'd14, 8'd229}: color_data = 12'h910;
			{9'd14, 8'd230}: color_data = 12'h200;
			{9'd14, 8'd231}: color_data = 12'h400;
			{9'd14, 8'd232}: color_data = 12'h900;
			{9'd14, 8'd233}: color_data = 12'ha00;
			{9'd14, 8'd234}: color_data = 12'h400;
			{9'd14, 8'd235}: color_data = 12'h310;
			{9'd14, 8'd236}: color_data = 12'hc30;
			{9'd14, 8'd237}: color_data = 12'hc20;
			{9'd14, 8'd238}: color_data = 12'h600;
			{9'd14, 8'd239}: color_data = 12'h000;
			{9'd15, 8'd16}: color_data = 12'h010;
			{9'd15, 8'd17}: color_data = 12'h780;
			{9'd15, 8'd18}: color_data = 12'hac0;
			{9'd15, 8'd19}: color_data = 12'hdea;
			{9'd15, 8'd20}: color_data = 12'hfff;
			{9'd15, 8'd21}: color_data = 12'hcd7;
			{9'd15, 8'd22}: color_data = 12'h8b0;
			{9'd15, 8'd23}: color_data = 12'h9b0;
			{9'd15, 8'd24}: color_data = 12'h9b0;
			{9'd15, 8'd25}: color_data = 12'h9b0;
			{9'd15, 8'd26}: color_data = 12'h9a0;
			{9'd15, 8'd27}: color_data = 12'h560;
			{9'd15, 8'd28}: color_data = 12'h120;
			{9'd15, 8'd29}: color_data = 12'h130;
			{9'd15, 8'd30}: color_data = 12'h240;
			{9'd15, 8'd31}: color_data = 12'h240;
			{9'd15, 8'd32}: color_data = 12'h140;
			{9'd15, 8'd33}: color_data = 12'h440;
			{9'd15, 8'd34}: color_data = 12'hc10;
			{9'd15, 8'd35}: color_data = 12'hf00;
			{9'd15, 8'd36}: color_data = 12'h720;
			{9'd15, 8'd37}: color_data = 12'h140;
			{9'd15, 8'd38}: color_data = 12'h920;
			{9'd15, 8'd39}: color_data = 12'hb10;
			{9'd15, 8'd40}: color_data = 12'h240;
			{9'd15, 8'd41}: color_data = 12'h530;
			{9'd15, 8'd42}: color_data = 12'he00;
			{9'd15, 8'd43}: color_data = 12'hd00;
			{9'd15, 8'd44}: color_data = 12'h430;
			{9'd15, 8'd45}: color_data = 12'h350;
			{9'd15, 8'd46}: color_data = 12'h790;
			{9'd15, 8'd47}: color_data = 12'h350;
			{9'd15, 8'd48}: color_data = 12'h030;
			{9'd15, 8'd49}: color_data = 12'h130;
			{9'd15, 8'd50}: color_data = 12'h020;
			{9'd15, 8'd51}: color_data = 12'h130;
			{9'd15, 8'd52}: color_data = 12'h240;
			{9'd15, 8'd53}: color_data = 12'h240;
			{9'd15, 8'd54}: color_data = 12'h240;
			{9'd15, 8'd55}: color_data = 12'h240;
			{9'd15, 8'd56}: color_data = 12'h240;
			{9'd15, 8'd57}: color_data = 12'h350;
			{9'd15, 8'd58}: color_data = 12'h560;
			{9'd15, 8'd59}: color_data = 12'h660;
			{9'd15, 8'd60}: color_data = 12'h760;
			{9'd15, 8'd61}: color_data = 12'h660;
			{9'd15, 8'd62}: color_data = 12'h220;
			{9'd15, 8'd63}: color_data = 12'h000;
			{9'd15, 8'd68}: color_data = 12'h047;
			{9'd15, 8'd69}: color_data = 12'h6df;
			{9'd15, 8'd70}: color_data = 12'hfff;
			{9'd15, 8'd71}: color_data = 12'hcbb;
			{9'd15, 8'd72}: color_data = 12'h323;
			{9'd15, 8'd73}: color_data = 12'h002;
			{9'd15, 8'd74}: color_data = 12'h000;
			{9'd15, 8'd75}: color_data = 12'h012;
			{9'd15, 8'd76}: color_data = 12'h08c;
			{9'd15, 8'd77}: color_data = 12'h034;
			{9'd15, 8'd128}: color_data = 12'h047;
			{9'd15, 8'd129}: color_data = 12'h6df;
			{9'd15, 8'd130}: color_data = 12'hfff;
			{9'd15, 8'd131}: color_data = 12'hcbb;
			{9'd15, 8'd132}: color_data = 12'h323;
			{9'd15, 8'd133}: color_data = 12'h002;
			{9'd15, 8'd134}: color_data = 12'h000;
			{9'd15, 8'd135}: color_data = 12'h012;
			{9'd15, 8'd136}: color_data = 12'h08c;
			{9'd15, 8'd137}: color_data = 12'h034;
			{9'd15, 8'd170}: color_data = 12'h000;
			{9'd15, 8'd171}: color_data = 12'h068;
			{9'd15, 8'd172}: color_data = 12'h8ef;
			{9'd15, 8'd173}: color_data = 12'hfff;
			{9'd15, 8'd174}: color_data = 12'haaa;
			{9'd15, 8'd175}: color_data = 12'h213;
			{9'd15, 8'd176}: color_data = 12'h002;
			{9'd15, 8'd178}: color_data = 12'h023;
			{9'd15, 8'd179}: color_data = 12'h08c;
			{9'd15, 8'd180}: color_data = 12'h023;
			{9'd15, 8'd204}: color_data = 12'h330;
			{9'd15, 8'd205}: color_data = 12'h790;
			{9'd15, 8'd206}: color_data = 12'h9b3;
			{9'd15, 8'd207}: color_data = 12'hcdd;
			{9'd15, 8'd208}: color_data = 12'hbca;
			{9'd15, 8'd209}: color_data = 12'h791;
			{9'd15, 8'd210}: color_data = 12'h790;
			{9'd15, 8'd211}: color_data = 12'h790;
			{9'd15, 8'd212}: color_data = 12'h790;
			{9'd15, 8'd213}: color_data = 12'h790;
			{9'd15, 8'd214}: color_data = 12'h790;
			{9'd15, 8'd215}: color_data = 12'h670;
			{9'd15, 8'd216}: color_data = 12'h230;
			{9'd15, 8'd217}: color_data = 12'h020;
			{9'd15, 8'd218}: color_data = 12'h130;
			{9'd15, 8'd219}: color_data = 12'h240;
			{9'd15, 8'd220}: color_data = 12'h550;
			{9'd15, 8'd221}: color_data = 12'h340;
			{9'd15, 8'd222}: color_data = 12'h200;
			{9'd15, 8'd223}: color_data = 12'h800;
			{9'd15, 8'd224}: color_data = 12'ha00;
			{9'd15, 8'd225}: color_data = 12'h800;
			{9'd15, 8'd226}: color_data = 12'h100;
			{9'd15, 8'd227}: color_data = 12'h100;
			{9'd15, 8'd228}: color_data = 12'h310;
			{9'd15, 8'd229}: color_data = 12'h200;
			{9'd15, 8'd230}: color_data = 12'h000;
			{9'd15, 8'd231}: color_data = 12'h500;
			{9'd15, 8'd232}: color_data = 12'ha00;
			{9'd15, 8'd233}: color_data = 12'ha00;
			{9'd15, 8'd234}: color_data = 12'h500;
			{9'd15, 8'd235}: color_data = 12'h000;
			{9'd15, 8'd236}: color_data = 12'h200;
			{9'd15, 8'd237}: color_data = 12'h300;
			{9'd15, 8'd238}: color_data = 12'h100;
			{9'd15, 8'd239}: color_data = 12'h000;
			{9'd16, 8'd16}: color_data = 12'h010;
			{9'd16, 8'd17}: color_data = 12'h780;
			{9'd16, 8'd18}: color_data = 12'hac0;
			{9'd16, 8'd19}: color_data = 12'hdea;
			{9'd16, 8'd20}: color_data = 12'hfff;
			{9'd16, 8'd21}: color_data = 12'hcd7;
			{9'd16, 8'd22}: color_data = 12'h9b0;
			{9'd16, 8'd23}: color_data = 12'h9b0;
			{9'd16, 8'd24}: color_data = 12'h9b0;
			{9'd16, 8'd25}: color_data = 12'h9a0;
			{9'd16, 8'd26}: color_data = 12'h660;
			{9'd16, 8'd27}: color_data = 12'h130;
			{9'd16, 8'd28}: color_data = 12'h130;
			{9'd16, 8'd29}: color_data = 12'h240;
			{9'd16, 8'd30}: color_data = 12'h140;
			{9'd16, 8'd31}: color_data = 12'h240;
			{9'd16, 8'd32}: color_data = 12'h450;
			{9'd16, 8'd33}: color_data = 12'h460;
			{9'd16, 8'd34}: color_data = 12'h750;
			{9'd16, 8'd35}: color_data = 12'he10;
			{9'd16, 8'd36}: color_data = 12'he00;
			{9'd16, 8'd37}: color_data = 12'hb10;
			{9'd16, 8'd38}: color_data = 12'hd00;
			{9'd16, 8'd39}: color_data = 12'he00;
			{9'd16, 8'd40}: color_data = 12'hb10;
			{9'd16, 8'd41}: color_data = 12'hd00;
			{9'd16, 8'd42}: color_data = 12'hf00;
			{9'd16, 8'd43}: color_data = 12'h940;
			{9'd16, 8'd44}: color_data = 12'h450;
			{9'd16, 8'd45}: color_data = 12'h560;
			{9'd16, 8'd46}: color_data = 12'h8a0;
			{9'd16, 8'd47}: color_data = 12'h460;
			{9'd16, 8'd48}: color_data = 12'h140;
			{9'd16, 8'd49}: color_data = 12'h240;
			{9'd16, 8'd50}: color_data = 12'h020;
			{9'd16, 8'd51}: color_data = 12'h240;
			{9'd16, 8'd52}: color_data = 12'h560;
			{9'd16, 8'd53}: color_data = 12'h550;
			{9'd16, 8'd54}: color_data = 12'h550;
			{9'd16, 8'd55}: color_data = 12'h550;
			{9'd16, 8'd56}: color_data = 12'h550;
			{9'd16, 8'd57}: color_data = 12'h560;
			{9'd16, 8'd58}: color_data = 12'h760;
			{9'd16, 8'd59}: color_data = 12'h770;
			{9'd16, 8'd60}: color_data = 12'h660;
			{9'd16, 8'd61}: color_data = 12'h220;
			{9'd16, 8'd62}: color_data = 12'h000;
			{9'd16, 8'd68}: color_data = 12'h047;
			{9'd16, 8'd69}: color_data = 12'h6ef;
			{9'd16, 8'd70}: color_data = 12'hddc;
			{9'd16, 8'd71}: color_data = 12'h434;
			{9'd16, 8'd72}: color_data = 12'h003;
			{9'd16, 8'd73}: color_data = 12'h005;
			{9'd16, 8'd74}: color_data = 12'h002;
			{9'd16, 8'd75}: color_data = 12'h012;
			{9'd16, 8'd76}: color_data = 12'h08c;
			{9'd16, 8'd77}: color_data = 12'h034;
			{9'd16, 8'd128}: color_data = 12'h047;
			{9'd16, 8'd129}: color_data = 12'h6ef;
			{9'd16, 8'd130}: color_data = 12'hddc;
			{9'd16, 8'd131}: color_data = 12'h434;
			{9'd16, 8'd132}: color_data = 12'h003;
			{9'd16, 8'd133}: color_data = 12'h005;
			{9'd16, 8'd134}: color_data = 12'h002;
			{9'd16, 8'd135}: color_data = 12'h012;
			{9'd16, 8'd136}: color_data = 12'h08c;
			{9'd16, 8'd137}: color_data = 12'h034;
			{9'd16, 8'd170}: color_data = 12'h000;
			{9'd16, 8'd171}: color_data = 12'h068;
			{9'd16, 8'd172}: color_data = 12'h8ff;
			{9'd16, 8'd173}: color_data = 12'hcbb;
			{9'd16, 8'd174}: color_data = 12'h323;
			{9'd16, 8'd175}: color_data = 12'h003;
			{9'd16, 8'd176}: color_data = 12'h005;
			{9'd16, 8'd177}: color_data = 12'h002;
			{9'd16, 8'd178}: color_data = 12'h023;
			{9'd16, 8'd179}: color_data = 12'h09c;
			{9'd16, 8'd180}: color_data = 12'h023;
			{9'd16, 8'd204}: color_data = 12'h340;
			{9'd16, 8'd205}: color_data = 12'h9c0;
			{9'd16, 8'd206}: color_data = 12'hcd4;
			{9'd16, 8'd207}: color_data = 12'hfff;
			{9'd16, 8'd208}: color_data = 12'hffd;
			{9'd16, 8'd209}: color_data = 12'hac1;
			{9'd16, 8'd210}: color_data = 12'h9b0;
			{9'd16, 8'd211}: color_data = 12'hac0;
			{9'd16, 8'd212}: color_data = 12'hac0;
			{9'd16, 8'd213}: color_data = 12'hac0;
			{9'd16, 8'd214}: color_data = 12'hac0;
			{9'd16, 8'd215}: color_data = 12'h890;
			{9'd16, 8'd216}: color_data = 12'h230;
			{9'd16, 8'd217}: color_data = 12'h030;
			{9'd16, 8'd218}: color_data = 12'h140;
			{9'd16, 8'd219}: color_data = 12'h450;
			{9'd16, 8'd220}: color_data = 12'h770;
			{9'd16, 8'd221}: color_data = 12'h440;
			{9'd16, 8'd222}: color_data = 12'h310;
			{9'd16, 8'd223}: color_data = 12'hc20;
			{9'd16, 8'd224}: color_data = 12'ha00;
			{9'd16, 8'd225}: color_data = 12'h800;
			{9'd16, 8'd226}: color_data = 12'h100;
			{9'd16, 8'd227}: color_data = 12'h300;
			{9'd16, 8'd228}: color_data = 12'h500;
			{9'd16, 8'd229}: color_data = 12'h500;
			{9'd16, 8'd230}: color_data = 12'h100;
			{9'd16, 8'd231}: color_data = 12'h710;
			{9'd16, 8'd232}: color_data = 12'hc10;
			{9'd16, 8'd233}: color_data = 12'h900;
			{9'd16, 8'd234}: color_data = 12'h500;
			{9'd16, 8'd235}: color_data = 12'h100;
			{9'd16, 8'd236}: color_data = 12'h500;
			{9'd16, 8'd237}: color_data = 12'h500;
			{9'd16, 8'd238}: color_data = 12'h400;
			{9'd16, 8'd239}: color_data = 12'h000;
			{9'd17, 8'd16}: color_data = 12'h010;
			{9'd17, 8'd17}: color_data = 12'h780;
			{9'd17, 8'd18}: color_data = 12'hac0;
			{9'd17, 8'd19}: color_data = 12'hdea;
			{9'd17, 8'd20}: color_data = 12'hfff;
			{9'd17, 8'd21}: color_data = 12'hcd7;
			{9'd17, 8'd22}: color_data = 12'h9b0;
			{9'd17, 8'd23}: color_data = 12'h9b0;
			{9'd17, 8'd24}: color_data = 12'h9b0;
			{9'd17, 8'd25}: color_data = 12'h8a0;
			{9'd17, 8'd26}: color_data = 12'h440;
			{9'd17, 8'd27}: color_data = 12'h020;
			{9'd17, 8'd28}: color_data = 12'h140;
			{9'd17, 8'd29}: color_data = 12'h240;
			{9'd17, 8'd30}: color_data = 12'h140;
			{9'd17, 8'd31}: color_data = 12'h350;
			{9'd17, 8'd32}: color_data = 12'h660;
			{9'd17, 8'd33}: color_data = 12'h770;
			{9'd17, 8'd34}: color_data = 12'h670;
			{9'd17, 8'd35}: color_data = 12'h950;
			{9'd17, 8'd36}: color_data = 12'hc30;
			{9'd17, 8'd37}: color_data = 12'hc30;
			{9'd17, 8'd38}: color_data = 12'hc30;
			{9'd17, 8'd39}: color_data = 12'hc30;
			{9'd17, 8'd40}: color_data = 12'hc30;
			{9'd17, 8'd41}: color_data = 12'hc30;
			{9'd17, 8'd42}: color_data = 12'ha40;
			{9'd17, 8'd43}: color_data = 12'h670;
			{9'd17, 8'd44}: color_data = 12'h670;
			{9'd17, 8'd45}: color_data = 12'h770;
			{9'd17, 8'd46}: color_data = 12'h8a0;
			{9'd17, 8'd47}: color_data = 12'h570;
			{9'd17, 8'd48}: color_data = 12'h450;
			{9'd17, 8'd49}: color_data = 12'h450;
			{9'd17, 8'd50}: color_data = 12'h130;
			{9'd17, 8'd51}: color_data = 12'h340;
			{9'd17, 8'd52}: color_data = 12'h770;
			{9'd17, 8'd53}: color_data = 12'h770;
			{9'd17, 8'd54}: color_data = 12'h770;
			{9'd17, 8'd55}: color_data = 12'h770;
			{9'd17, 8'd56}: color_data = 12'h770;
			{9'd17, 8'd57}: color_data = 12'h660;
			{9'd17, 8'd58}: color_data = 12'h330;
			{9'd17, 8'd59}: color_data = 12'h330;
			{9'd17, 8'd60}: color_data = 12'h220;
			{9'd17, 8'd61}: color_data = 12'h000;
			{9'd17, 8'd68}: color_data = 12'h057;
			{9'd17, 8'd69}: color_data = 12'h3bd;
			{9'd17, 8'd70}: color_data = 12'h555;
			{9'd17, 8'd71}: color_data = 12'h002;
			{9'd17, 8'd72}: color_data = 12'h005;
			{9'd17, 8'd73}: color_data = 12'h005;
			{9'd17, 8'd74}: color_data = 12'h004;
			{9'd17, 8'd75}: color_data = 12'h025;
			{9'd17, 8'd76}: color_data = 12'h09c;
			{9'd17, 8'd77}: color_data = 12'h034;
			{9'd17, 8'd128}: color_data = 12'h057;
			{9'd17, 8'd129}: color_data = 12'h3bd;
			{9'd17, 8'd130}: color_data = 12'h555;
			{9'd17, 8'd131}: color_data = 12'h002;
			{9'd17, 8'd132}: color_data = 12'h005;
			{9'd17, 8'd133}: color_data = 12'h005;
			{9'd17, 8'd134}: color_data = 12'h004;
			{9'd17, 8'd135}: color_data = 12'h024;
			{9'd17, 8'd136}: color_data = 12'h09c;
			{9'd17, 8'd137}: color_data = 12'h034;
			{9'd17, 8'd170}: color_data = 12'h000;
			{9'd17, 8'd171}: color_data = 12'h079;
			{9'd17, 8'd172}: color_data = 12'h4bd;
			{9'd17, 8'd173}: color_data = 12'h444;
			{9'd17, 8'd174}: color_data = 12'h002;
			{9'd17, 8'd175}: color_data = 12'h005;
			{9'd17, 8'd176}: color_data = 12'h005;
			{9'd17, 8'd177}: color_data = 12'h004;
			{9'd17, 8'd178}: color_data = 12'h036;
			{9'd17, 8'd179}: color_data = 12'h09c;
			{9'd17, 8'd180}: color_data = 12'h023;
			{9'd17, 8'd204}: color_data = 12'h340;
			{9'd17, 8'd205}: color_data = 12'h9b0;
			{9'd17, 8'd206}: color_data = 12'hbc4;
			{9'd17, 8'd207}: color_data = 12'hfff;
			{9'd17, 8'd208}: color_data = 12'hefd;
			{9'd17, 8'd209}: color_data = 12'h9b1;
			{9'd17, 8'd210}: color_data = 12'h9b0;
			{9'd17, 8'd211}: color_data = 12'h9b0;
			{9'd17, 8'd212}: color_data = 12'h9b0;
			{9'd17, 8'd213}: color_data = 12'h9b0;
			{9'd17, 8'd214}: color_data = 12'h9b0;
			{9'd17, 8'd215}: color_data = 12'h780;
			{9'd17, 8'd216}: color_data = 12'h230;
			{9'd17, 8'd217}: color_data = 12'h020;
			{9'd17, 8'd218}: color_data = 12'h140;
			{9'd17, 8'd219}: color_data = 12'h350;
			{9'd17, 8'd220}: color_data = 12'h770;
			{9'd17, 8'd221}: color_data = 12'h340;
			{9'd17, 8'd222}: color_data = 12'h410;
			{9'd17, 8'd223}: color_data = 12'hd30;
			{9'd17, 8'd224}: color_data = 12'hb00;
			{9'd17, 8'd225}: color_data = 12'h700;
			{9'd17, 8'd226}: color_data = 12'h200;
			{9'd17, 8'd227}: color_data = 12'h700;
			{9'd17, 8'd228}: color_data = 12'hb00;
			{9'd17, 8'd229}: color_data = 12'ha00;
			{9'd17, 8'd230}: color_data = 12'h300;
			{9'd17, 8'd231}: color_data = 12'h820;
			{9'd17, 8'd232}: color_data = 12'hd20;
			{9'd17, 8'd233}: color_data = 12'h900;
			{9'd17, 8'd234}: color_data = 12'h500;
			{9'd17, 8'd235}: color_data = 12'h300;
			{9'd17, 8'd236}: color_data = 12'h900;
			{9'd17, 8'd237}: color_data = 12'hb00;
			{9'd17, 8'd238}: color_data = 12'h800;
			{9'd17, 8'd239}: color_data = 12'h100;
			{9'd18, 8'd16}: color_data = 12'h010;
			{9'd18, 8'd17}: color_data = 12'h780;
			{9'd18, 8'd18}: color_data = 12'hac0;
			{9'd18, 8'd19}: color_data = 12'hdea;
			{9'd18, 8'd20}: color_data = 12'hfff;
			{9'd18, 8'd21}: color_data = 12'hcd7;
			{9'd18, 8'd22}: color_data = 12'h9b0;
			{9'd18, 8'd23}: color_data = 12'h9b0;
			{9'd18, 8'd24}: color_data = 12'h9b0;
			{9'd18, 8'd25}: color_data = 12'h8a0;
			{9'd18, 8'd26}: color_data = 12'h450;
			{9'd18, 8'd27}: color_data = 12'h020;
			{9'd18, 8'd28}: color_data = 12'h140;
			{9'd18, 8'd29}: color_data = 12'h240;
			{9'd18, 8'd30}: color_data = 12'h350;
			{9'd18, 8'd31}: color_data = 12'h660;
			{9'd18, 8'd32}: color_data = 12'h760;
			{9'd18, 8'd33}: color_data = 12'h550;
			{9'd18, 8'd34}: color_data = 12'h440;
			{9'd18, 8'd35}: color_data = 12'h440;
			{9'd18, 8'd36}: color_data = 12'h440;
			{9'd18, 8'd37}: color_data = 12'h440;
			{9'd18, 8'd38}: color_data = 12'h440;
			{9'd18, 8'd39}: color_data = 12'h440;
			{9'd18, 8'd40}: color_data = 12'h440;
			{9'd18, 8'd41}: color_data = 12'h440;
			{9'd18, 8'd42}: color_data = 12'h440;
			{9'd18, 8'd43}: color_data = 12'h440;
			{9'd18, 8'd44}: color_data = 12'h440;
			{9'd18, 8'd45}: color_data = 12'h550;
			{9'd18, 8'd46}: color_data = 12'h8a0;
			{9'd18, 8'd47}: color_data = 12'h880;
			{9'd18, 8'd48}: color_data = 12'h760;
			{9'd18, 8'd49}: color_data = 12'h770;
			{9'd18, 8'd50}: color_data = 12'h230;
			{9'd18, 8'd51}: color_data = 12'h220;
			{9'd18, 8'd52}: color_data = 12'h440;
			{9'd18, 8'd53}: color_data = 12'h440;
			{9'd18, 8'd54}: color_data = 12'h440;
			{9'd18, 8'd55}: color_data = 12'h440;
			{9'd18, 8'd56}: color_data = 12'h440;
			{9'd18, 8'd57}: color_data = 12'h330;
			{9'd18, 8'd58}: color_data = 12'h000;
			{9'd18, 8'd60}: color_data = 12'h000;
			{9'd18, 8'd68}: color_data = 12'h035;
			{9'd18, 8'd69}: color_data = 12'h047;
			{9'd18, 8'd70}: color_data = 12'h001;
			{9'd18, 8'd71}: color_data = 12'h004;
			{9'd18, 8'd72}: color_data = 12'h004;
			{9'd18, 8'd73}: color_data = 12'h004;
			{9'd18, 8'd74}: color_data = 12'h004;
			{9'd18, 8'd75}: color_data = 12'h015;
			{9'd18, 8'd76}: color_data = 12'h059;
			{9'd18, 8'd77}: color_data = 12'h023;
			{9'd18, 8'd128}: color_data = 12'h035;
			{9'd18, 8'd129}: color_data = 12'h047;
			{9'd18, 8'd130}: color_data = 12'h001;
			{9'd18, 8'd131}: color_data = 12'h004;
			{9'd18, 8'd132}: color_data = 12'h004;
			{9'd18, 8'd133}: color_data = 12'h004;
			{9'd18, 8'd134}: color_data = 12'h004;
			{9'd18, 8'd135}: color_data = 12'h015;
			{9'd18, 8'd136}: color_data = 12'h059;
			{9'd18, 8'd137}: color_data = 12'h023;
			{9'd18, 8'd170}: color_data = 12'h000;
			{9'd18, 8'd171}: color_data = 12'h047;
			{9'd18, 8'd172}: color_data = 12'h036;
			{9'd18, 8'd173}: color_data = 12'h001;
			{9'd18, 8'd174}: color_data = 12'h004;
			{9'd18, 8'd175}: color_data = 12'h004;
			{9'd18, 8'd176}: color_data = 12'h004;
			{9'd18, 8'd177}: color_data = 12'h004;
			{9'd18, 8'd178}: color_data = 12'h016;
			{9'd18, 8'd179}: color_data = 12'h059;
			{9'd18, 8'd180}: color_data = 12'h012;
			{9'd18, 8'd204}: color_data = 12'h340;
			{9'd18, 8'd205}: color_data = 12'had1;
			{9'd18, 8'd206}: color_data = 12'hdf9;
			{9'd18, 8'd207}: color_data = 12'hfff;
			{9'd18, 8'd208}: color_data = 12'hffe;
			{9'd18, 8'd209}: color_data = 12'hce6;
			{9'd18, 8'd210}: color_data = 12'hac0;
			{9'd18, 8'd211}: color_data = 12'h9c0;
			{9'd18, 8'd212}: color_data = 12'hac0;
			{9'd18, 8'd213}: color_data = 12'hac0;
			{9'd18, 8'd214}: color_data = 12'hac0;
			{9'd18, 8'd215}: color_data = 12'h890;
			{9'd18, 8'd216}: color_data = 12'h230;
			{9'd18, 8'd217}: color_data = 12'h030;
			{9'd18, 8'd218}: color_data = 12'h140;
			{9'd18, 8'd219}: color_data = 12'h450;
			{9'd18, 8'd220}: color_data = 12'h770;
			{9'd18, 8'd221}: color_data = 12'h440;
			{9'd18, 8'd222}: color_data = 12'h410;
			{9'd18, 8'd223}: color_data = 12'he30;
			{9'd18, 8'd224}: color_data = 12'hd20;
			{9'd18, 8'd225}: color_data = 12'h800;
			{9'd18, 8'd226}: color_data = 12'h200;
			{9'd18, 8'd227}: color_data = 12'h600;
			{9'd18, 8'd228}: color_data = 12'ha00;
			{9'd18, 8'd229}: color_data = 12'h900;
			{9'd18, 8'd230}: color_data = 12'h300;
			{9'd18, 8'd231}: color_data = 12'h820;
			{9'd18, 8'd232}: color_data = 12'hf30;
			{9'd18, 8'd233}: color_data = 12'hc00;
			{9'd18, 8'd234}: color_data = 12'h500;
			{9'd18, 8'd235}: color_data = 12'h200;
			{9'd18, 8'd236}: color_data = 12'h900;
			{9'd18, 8'd237}: color_data = 12'ha00;
			{9'd18, 8'd238}: color_data = 12'h700;
			{9'd18, 8'd239}: color_data = 12'h100;
			{9'd19, 8'd16}: color_data = 12'h010;
			{9'd19, 8'd17}: color_data = 12'h780;
			{9'd19, 8'd18}: color_data = 12'hac0;
			{9'd19, 8'd19}: color_data = 12'hdea;
			{9'd19, 8'd20}: color_data = 12'hfff;
			{9'd19, 8'd21}: color_data = 12'hcd7;
			{9'd19, 8'd22}: color_data = 12'h9b0;
			{9'd19, 8'd23}: color_data = 12'h9b0;
			{9'd19, 8'd24}: color_data = 12'h9b0;
			{9'd19, 8'd25}: color_data = 12'h8a0;
			{9'd19, 8'd26}: color_data = 12'h450;
			{9'd19, 8'd27}: color_data = 12'h020;
			{9'd19, 8'd28}: color_data = 12'h140;
			{9'd19, 8'd29}: color_data = 12'h240;
			{9'd19, 8'd30}: color_data = 12'h560;
			{9'd19, 8'd31}: color_data = 12'h660;
			{9'd19, 8'd32}: color_data = 12'h550;
			{9'd19, 8'd33}: color_data = 12'h110;
			{9'd19, 8'd34}: color_data = 12'h000;
			{9'd19, 8'd35}: color_data = 12'h000;
			{9'd19, 8'd36}: color_data = 12'h000;
			{9'd19, 8'd37}: color_data = 12'h000;
			{9'd19, 8'd38}: color_data = 12'h000;
			{9'd19, 8'd39}: color_data = 12'h000;
			{9'd19, 8'd40}: color_data = 12'h000;
			{9'd19, 8'd41}: color_data = 12'h000;
			{9'd19, 8'd42}: color_data = 12'h000;
			{9'd19, 8'd43}: color_data = 12'h000;
			{9'd19, 8'd44}: color_data = 12'h000;
			{9'd19, 8'd45}: color_data = 12'h110;
			{9'd19, 8'd46}: color_data = 12'h670;
			{9'd19, 8'd47}: color_data = 12'h670;
			{9'd19, 8'd48}: color_data = 12'h550;
			{9'd19, 8'd49}: color_data = 12'h550;
			{9'd19, 8'd50}: color_data = 12'h220;
			{9'd19, 8'd51}: color_data = 12'h000;
			{9'd19, 8'd52}: color_data = 12'h000;
			{9'd19, 8'd53}: color_data = 12'h000;
			{9'd19, 8'd54}: color_data = 12'h000;
			{9'd19, 8'd55}: color_data = 12'h000;
			{9'd19, 8'd56}: color_data = 12'h000;
			{9'd19, 8'd57}: color_data = 12'h000;
			{9'd19, 8'd68}: color_data = 12'h013;
			{9'd19, 8'd69}: color_data = 12'h027;
			{9'd19, 8'd70}: color_data = 12'h016;
			{9'd19, 8'd71}: color_data = 12'h027;
			{9'd19, 8'd72}: color_data = 12'h027;
			{9'd19, 8'd73}: color_data = 12'h027;
			{9'd19, 8'd74}: color_data = 12'h027;
			{9'd19, 8'd75}: color_data = 12'h028;
			{9'd19, 8'd76}: color_data = 12'h027;
			{9'd19, 8'd77}: color_data = 12'h001;
			{9'd19, 8'd128}: color_data = 12'h013;
			{9'd19, 8'd129}: color_data = 12'h027;
			{9'd19, 8'd130}: color_data = 12'h016;
			{9'd19, 8'd131}: color_data = 12'h027;
			{9'd19, 8'd132}: color_data = 12'h027;
			{9'd19, 8'd133}: color_data = 12'h027;
			{9'd19, 8'd134}: color_data = 12'h027;
			{9'd19, 8'd135}: color_data = 12'h028;
			{9'd19, 8'd136}: color_data = 12'h027;
			{9'd19, 8'd137}: color_data = 12'h001;
			{9'd19, 8'd170}: color_data = 12'h000;
			{9'd19, 8'd171}: color_data = 12'h014;
			{9'd19, 8'd172}: color_data = 12'h027;
			{9'd19, 8'd173}: color_data = 12'h016;
			{9'd19, 8'd174}: color_data = 12'h027;
			{9'd19, 8'd175}: color_data = 12'h027;
			{9'd19, 8'd176}: color_data = 12'h027;
			{9'd19, 8'd177}: color_data = 12'h027;
			{9'd19, 8'd178}: color_data = 12'h028;
			{9'd19, 8'd179}: color_data = 12'h026;
			{9'd19, 8'd180}: color_data = 12'h001;
			{9'd19, 8'd204}: color_data = 12'h230;
			{9'd19, 8'd205}: color_data = 12'h9b4;
			{9'd19, 8'd206}: color_data = 12'hddc;
			{9'd19, 8'd207}: color_data = 12'hddd;
			{9'd19, 8'd208}: color_data = 12'hddd;
			{9'd19, 8'd209}: color_data = 12'hccb;
			{9'd19, 8'd210}: color_data = 12'h8a1;
			{9'd19, 8'd211}: color_data = 12'h790;
			{9'd19, 8'd212}: color_data = 12'h790;
			{9'd19, 8'd213}: color_data = 12'h790;
			{9'd19, 8'd214}: color_data = 12'h890;
			{9'd19, 8'd215}: color_data = 12'h670;
			{9'd19, 8'd216}: color_data = 12'h230;
			{9'd19, 8'd217}: color_data = 12'h020;
			{9'd19, 8'd218}: color_data = 12'h130;
			{9'd19, 8'd219}: color_data = 12'h340;
			{9'd19, 8'd220}: color_data = 12'h550;
			{9'd19, 8'd221}: color_data = 12'h330;
			{9'd19, 8'd222}: color_data = 12'h200;
			{9'd19, 8'd223}: color_data = 12'hb30;
			{9'd19, 8'd224}: color_data = 12'hc30;
			{9'd19, 8'd225}: color_data = 12'h600;
			{9'd19, 8'd226}: color_data = 12'h100;
			{9'd19, 8'd227}: color_data = 12'h600;
			{9'd19, 8'd228}: color_data = 12'ha00;
			{9'd19, 8'd229}: color_data = 12'h900;
			{9'd19, 8'd230}: color_data = 12'h300;
			{9'd19, 8'd231}: color_data = 12'h620;
			{9'd19, 8'd232}: color_data = 12'hd40;
			{9'd19, 8'd233}: color_data = 12'ha20;
			{9'd19, 8'd234}: color_data = 12'h300;
			{9'd19, 8'd235}: color_data = 12'h200;
			{9'd19, 8'd236}: color_data = 12'h900;
			{9'd19, 8'd237}: color_data = 12'ha00;
			{9'd19, 8'd238}: color_data = 12'h700;
			{9'd19, 8'd239}: color_data = 12'h100;
			{9'd20, 8'd16}: color_data = 12'h010;
			{9'd20, 8'd17}: color_data = 12'h780;
			{9'd20, 8'd18}: color_data = 12'hac0;
			{9'd20, 8'd19}: color_data = 12'hdea;
			{9'd20, 8'd20}: color_data = 12'hfff;
			{9'd20, 8'd21}: color_data = 12'hcd7;
			{9'd20, 8'd22}: color_data = 12'h9b0;
			{9'd20, 8'd23}: color_data = 12'h9b0;
			{9'd20, 8'd24}: color_data = 12'h9b0;
			{9'd20, 8'd25}: color_data = 12'h8a0;
			{9'd20, 8'd26}: color_data = 12'h450;
			{9'd20, 8'd27}: color_data = 12'h020;
			{9'd20, 8'd28}: color_data = 12'h140;
			{9'd20, 8'd29}: color_data = 12'h240;
			{9'd20, 8'd30}: color_data = 12'h660;
			{9'd20, 8'd31}: color_data = 12'h660;
			{9'd20, 8'd32}: color_data = 12'h220;
			{9'd20, 8'd33}: color_data = 12'h000;
			{9'd20, 8'd45}: color_data = 12'h000;
			{9'd20, 8'd46}: color_data = 12'h110;
			{9'd20, 8'd47}: color_data = 12'h110;
			{9'd20, 8'd48}: color_data = 12'h110;
			{9'd20, 8'd49}: color_data = 12'h110;
			{9'd20, 8'd50}: color_data = 12'h000;
			{9'd20, 8'd68}: color_data = 12'h035;
			{9'd20, 8'd69}: color_data = 12'h09e;
			{9'd20, 8'd70}: color_data = 12'h09e;
			{9'd20, 8'd71}: color_data = 12'h09e;
			{9'd20, 8'd72}: color_data = 12'h09e;
			{9'd20, 8'd73}: color_data = 12'h09e;
			{9'd20, 8'd74}: color_data = 12'h09e;
			{9'd20, 8'd75}: color_data = 12'h09e;
			{9'd20, 8'd76}: color_data = 12'h08c;
			{9'd20, 8'd77}: color_data = 12'h023;
			{9'd20, 8'd128}: color_data = 12'h035;
			{9'd20, 8'd129}: color_data = 12'h09e;
			{9'd20, 8'd130}: color_data = 12'h09e;
			{9'd20, 8'd131}: color_data = 12'h09e;
			{9'd20, 8'd132}: color_data = 12'h09e;
			{9'd20, 8'd133}: color_data = 12'h09e;
			{9'd20, 8'd134}: color_data = 12'h09e;
			{9'd20, 8'd135}: color_data = 12'h09e;
			{9'd20, 8'd136}: color_data = 12'h08c;
			{9'd20, 8'd137}: color_data = 12'h023;
			{9'd20, 8'd170}: color_data = 12'h000;
			{9'd20, 8'd171}: color_data = 12'h057;
			{9'd20, 8'd172}: color_data = 12'h0ae;
			{9'd20, 8'd173}: color_data = 12'h09e;
			{9'd20, 8'd174}: color_data = 12'h09e;
			{9'd20, 8'd175}: color_data = 12'h09e;
			{9'd20, 8'd176}: color_data = 12'h09e;
			{9'd20, 8'd177}: color_data = 12'h09e;
			{9'd20, 8'd178}: color_data = 12'h09e;
			{9'd20, 8'd179}: color_data = 12'h07b;
			{9'd20, 8'd180}: color_data = 12'h012;
			{9'd20, 8'd204}: color_data = 12'h000;
			{9'd20, 8'd205}: color_data = 12'h221;
			{9'd20, 8'd206}: color_data = 12'h333;
			{9'd20, 8'd207}: color_data = 12'h222;
			{9'd20, 8'd208}: color_data = 12'h223;
			{9'd20, 8'd209}: color_data = 12'h223;
			{9'd20, 8'd210}: color_data = 12'h120;
			{9'd20, 8'd211}: color_data = 12'h110;
			{9'd20, 8'd212}: color_data = 12'h120;
			{9'd20, 8'd213}: color_data = 12'h120;
			{9'd20, 8'd214}: color_data = 12'h120;
			{9'd20, 8'd215}: color_data = 12'h110;
			{9'd20, 8'd216}: color_data = 12'h000;
			{9'd20, 8'd217}: color_data = 12'h000;
			{9'd20, 8'd218}: color_data = 12'h000;
			{9'd20, 8'd219}: color_data = 12'h000;
			{9'd20, 8'd220}: color_data = 12'h110;
			{9'd20, 8'd221}: color_data = 12'h000;
			{9'd20, 8'd222}: color_data = 12'h000;
			{9'd20, 8'd223}: color_data = 12'h200;
			{9'd20, 8'd224}: color_data = 12'h300;
			{9'd20, 8'd225}: color_data = 12'h100;
			{9'd20, 8'd226}: color_data = 12'h000;
			{9'd20, 8'd227}: color_data = 12'h700;
			{9'd20, 8'd228}: color_data = 12'ha00;
			{9'd20, 8'd229}: color_data = 12'h900;
			{9'd20, 8'd230}: color_data = 12'h300;
			{9'd20, 8'd231}: color_data = 12'h100;
			{9'd20, 8'd232}: color_data = 12'h310;
			{9'd20, 8'd233}: color_data = 12'h200;
			{9'd20, 8'd234}: color_data = 12'h000;
			{9'd20, 8'd235}: color_data = 12'h300;
			{9'd20, 8'd236}: color_data = 12'h900;
			{9'd20, 8'd237}: color_data = 12'ha00;
			{9'd20, 8'd238}: color_data = 12'h700;
			{9'd20, 8'd239}: color_data = 12'h100;
			{9'd21, 8'd16}: color_data = 12'h010;
			{9'd21, 8'd17}: color_data = 12'h780;
			{9'd21, 8'd18}: color_data = 12'hac0;
			{9'd21, 8'd19}: color_data = 12'hdea;
			{9'd21, 8'd20}: color_data = 12'hfff;
			{9'd21, 8'd21}: color_data = 12'hcd7;
			{9'd21, 8'd22}: color_data = 12'h9b0;
			{9'd21, 8'd23}: color_data = 12'h9b0;
			{9'd21, 8'd24}: color_data = 12'h9b0;
			{9'd21, 8'd25}: color_data = 12'h8a0;
			{9'd21, 8'd26}: color_data = 12'h450;
			{9'd21, 8'd27}: color_data = 12'h020;
			{9'd21, 8'd28}: color_data = 12'h140;
			{9'd21, 8'd29}: color_data = 12'h240;
			{9'd21, 8'd30}: color_data = 12'h660;
			{9'd21, 8'd31}: color_data = 12'h660;
			{9'd21, 8'd32}: color_data = 12'h110;
			{9'd21, 8'd68}: color_data = 12'h057;
			{9'd21, 8'd69}: color_data = 12'h4ef;
			{9'd21, 8'd70}: color_data = 12'h7ef;
			{9'd21, 8'd71}: color_data = 12'h0cf;
			{9'd21, 8'd72}: color_data = 12'h0cf;
			{9'd21, 8'd73}: color_data = 12'h0df;
			{9'd21, 8'd74}: color_data = 12'h0bd;
			{9'd21, 8'd75}: color_data = 12'h068;
			{9'd21, 8'd76}: color_data = 12'h09c;
			{9'd21, 8'd77}: color_data = 12'h034;
			{9'd21, 8'd128}: color_data = 12'h057;
			{9'd21, 8'd129}: color_data = 12'h4ef;
			{9'd21, 8'd130}: color_data = 12'h7ef;
			{9'd21, 8'd131}: color_data = 12'h0cf;
			{9'd21, 8'd132}: color_data = 12'h0cf;
			{9'd21, 8'd133}: color_data = 12'h0df;
			{9'd21, 8'd134}: color_data = 12'h0bd;
			{9'd21, 8'd135}: color_data = 12'h068;
			{9'd21, 8'd136}: color_data = 12'h09c;
			{9'd21, 8'd137}: color_data = 12'h034;
			{9'd21, 8'd170}: color_data = 12'h000;
			{9'd21, 8'd171}: color_data = 12'h069;
			{9'd21, 8'd172}: color_data = 12'h6ef;
			{9'd21, 8'd173}: color_data = 12'h6ef;
			{9'd21, 8'd174}: color_data = 12'h0cf;
			{9'd21, 8'd175}: color_data = 12'h0cf;
			{9'd21, 8'd176}: color_data = 12'h0df;
			{9'd21, 8'd177}: color_data = 12'h0ac;
			{9'd21, 8'd178}: color_data = 12'h079;
			{9'd21, 8'd179}: color_data = 12'h09c;
			{9'd21, 8'd180}: color_data = 12'h023;
			{9'd21, 8'd222}: color_data = 12'h100;
			{9'd21, 8'd223}: color_data = 12'h400;
			{9'd21, 8'd224}: color_data = 12'h500;
			{9'd21, 8'd225}: color_data = 12'h400;
			{9'd21, 8'd226}: color_data = 12'h200;
			{9'd21, 8'd227}: color_data = 12'ha20;
			{9'd21, 8'd228}: color_data = 12'hb10;
			{9'd21, 8'd229}: color_data = 12'h900;
			{9'd21, 8'd230}: color_data = 12'h300;
			{9'd21, 8'd231}: color_data = 12'h200;
			{9'd21, 8'd232}: color_data = 12'h500;
			{9'd21, 8'd233}: color_data = 12'h500;
			{9'd21, 8'd234}: color_data = 12'h200;
			{9'd21, 8'd235}: color_data = 12'h410;
			{9'd21, 8'd236}: color_data = 12'hc20;
			{9'd21, 8'd237}: color_data = 12'ha00;
			{9'd21, 8'd238}: color_data = 12'h700;
			{9'd21, 8'd239}: color_data = 12'h100;
			{9'd22, 8'd16}: color_data = 12'h010;
			{9'd22, 8'd17}: color_data = 12'h780;
			{9'd22, 8'd18}: color_data = 12'hac0;
			{9'd22, 8'd19}: color_data = 12'hdea;
			{9'd22, 8'd20}: color_data = 12'hfff;
			{9'd22, 8'd21}: color_data = 12'hcd7;
			{9'd22, 8'd22}: color_data = 12'h9b0;
			{9'd22, 8'd23}: color_data = 12'h9b0;
			{9'd22, 8'd24}: color_data = 12'h9b0;
			{9'd22, 8'd25}: color_data = 12'h8a0;
			{9'd22, 8'd26}: color_data = 12'h450;
			{9'd22, 8'd27}: color_data = 12'h020;
			{9'd22, 8'd28}: color_data = 12'h140;
			{9'd22, 8'd29}: color_data = 12'h240;
			{9'd22, 8'd30}: color_data = 12'h660;
			{9'd22, 8'd31}: color_data = 12'h660;
			{9'd22, 8'd32}: color_data = 12'h110;
			{9'd22, 8'd68}: color_data = 12'h047;
			{9'd22, 8'd69}: color_data = 12'h6df;
			{9'd22, 8'd70}: color_data = 12'heff;
			{9'd22, 8'd71}: color_data = 12'h6df;
			{9'd22, 8'd72}: color_data = 12'h0bf;
			{9'd22, 8'd73}: color_data = 12'h0bf;
			{9'd22, 8'd74}: color_data = 12'h056;
			{9'd22, 8'd75}: color_data = 12'h012;
			{9'd22, 8'd76}: color_data = 12'h08b;
			{9'd22, 8'd77}: color_data = 12'h034;
			{9'd22, 8'd128}: color_data = 12'h047;
			{9'd22, 8'd129}: color_data = 12'h6df;
			{9'd22, 8'd130}: color_data = 12'heff;
			{9'd22, 8'd131}: color_data = 12'h6df;
			{9'd22, 8'd132}: color_data = 12'h0bf;
			{9'd22, 8'd133}: color_data = 12'h0bf;
			{9'd22, 8'd134}: color_data = 12'h056;
			{9'd22, 8'd135}: color_data = 12'h012;
			{9'd22, 8'd136}: color_data = 12'h08b;
			{9'd22, 8'd137}: color_data = 12'h034;
			{9'd22, 8'd170}: color_data = 12'h000;
			{9'd22, 8'd171}: color_data = 12'h068;
			{9'd22, 8'd172}: color_data = 12'h8ef;
			{9'd22, 8'd173}: color_data = 12'hdff;
			{9'd22, 8'd174}: color_data = 12'h4cf;
			{9'd22, 8'd175}: color_data = 12'h0cf;
			{9'd22, 8'd176}: color_data = 12'h0ae;
			{9'd22, 8'd177}: color_data = 12'h035;
			{9'd22, 8'd178}: color_data = 12'h023;
			{9'd22, 8'd179}: color_data = 12'h08c;
			{9'd22, 8'd180}: color_data = 12'h023;
			{9'd22, 8'd222}: color_data = 12'h200;
			{9'd22, 8'd223}: color_data = 12'h900;
			{9'd22, 8'd224}: color_data = 12'hb00;
			{9'd22, 8'd225}: color_data = 12'h800;
			{9'd22, 8'd226}: color_data = 12'h200;
			{9'd22, 8'd227}: color_data = 12'hb30;
			{9'd22, 8'd228}: color_data = 12'hc10;
			{9'd22, 8'd229}: color_data = 12'h800;
			{9'd22, 8'd230}: color_data = 12'h300;
			{9'd22, 8'd231}: color_data = 12'h400;
			{9'd22, 8'd232}: color_data = 12'ha00;
			{9'd22, 8'd233}: color_data = 12'ha00;
			{9'd22, 8'd234}: color_data = 12'h500;
			{9'd22, 8'd235}: color_data = 12'h510;
			{9'd22, 8'd236}: color_data = 12'hd30;
			{9'd22, 8'd237}: color_data = 12'ha00;
			{9'd22, 8'd238}: color_data = 12'h700;
			{9'd22, 8'd239}: color_data = 12'h100;
			{9'd23, 8'd16}: color_data = 12'h010;
			{9'd23, 8'd17}: color_data = 12'h780;
			{9'd23, 8'd18}: color_data = 12'hac0;
			{9'd23, 8'd19}: color_data = 12'hdea;
			{9'd23, 8'd20}: color_data = 12'hfff;
			{9'd23, 8'd21}: color_data = 12'hcd7;
			{9'd23, 8'd22}: color_data = 12'h9b0;
			{9'd23, 8'd23}: color_data = 12'h9b0;
			{9'd23, 8'd24}: color_data = 12'h9b0;
			{9'd23, 8'd25}: color_data = 12'h8a0;
			{9'd23, 8'd26}: color_data = 12'h450;
			{9'd23, 8'd27}: color_data = 12'h020;
			{9'd23, 8'd28}: color_data = 12'h140;
			{9'd23, 8'd29}: color_data = 12'h240;
			{9'd23, 8'd30}: color_data = 12'h660;
			{9'd23, 8'd31}: color_data = 12'h660;
			{9'd23, 8'd32}: color_data = 12'h110;
			{9'd23, 8'd68}: color_data = 12'h047;
			{9'd23, 8'd69}: color_data = 12'h6df;
			{9'd23, 8'd70}: color_data = 12'hfff;
			{9'd23, 8'd71}: color_data = 12'hdff;
			{9'd23, 8'd72}: color_data = 12'h5df;
			{9'd23, 8'd73}: color_data = 12'h068;
			{9'd23, 8'd74}: color_data = 12'h000;
			{9'd23, 8'd75}: color_data = 12'h012;
			{9'd23, 8'd76}: color_data = 12'h08c;
			{9'd23, 8'd77}: color_data = 12'h034;
			{9'd23, 8'd128}: color_data = 12'h047;
			{9'd23, 8'd129}: color_data = 12'h6df;
			{9'd23, 8'd130}: color_data = 12'hfff;
			{9'd23, 8'd131}: color_data = 12'hdff;
			{9'd23, 8'd132}: color_data = 12'h5df;
			{9'd23, 8'd133}: color_data = 12'h068;
			{9'd23, 8'd134}: color_data = 12'h000;
			{9'd23, 8'd135}: color_data = 12'h012;
			{9'd23, 8'd136}: color_data = 12'h08c;
			{9'd23, 8'd137}: color_data = 12'h034;
			{9'd23, 8'd170}: color_data = 12'h000;
			{9'd23, 8'd171}: color_data = 12'h068;
			{9'd23, 8'd172}: color_data = 12'h8ef;
			{9'd23, 8'd173}: color_data = 12'hfff;
			{9'd23, 8'd174}: color_data = 12'hcff;
			{9'd23, 8'd175}: color_data = 12'h4ce;
			{9'd23, 8'd176}: color_data = 12'h057;
			{9'd23, 8'd177}: color_data = 12'h000;
			{9'd23, 8'd178}: color_data = 12'h023;
			{9'd23, 8'd179}: color_data = 12'h08c;
			{9'd23, 8'd180}: color_data = 12'h023;
			{9'd23, 8'd222}: color_data = 12'h200;
			{9'd23, 8'd223}: color_data = 12'h900;
			{9'd23, 8'd224}: color_data = 12'ha00;
			{9'd23, 8'd225}: color_data = 12'h700;
			{9'd23, 8'd226}: color_data = 12'h200;
			{9'd23, 8'd227}: color_data = 12'hb30;
			{9'd23, 8'd228}: color_data = 12'he20;
			{9'd23, 8'd229}: color_data = 12'ha00;
			{9'd23, 8'd230}: color_data = 12'h300;
			{9'd23, 8'd231}: color_data = 12'h400;
			{9'd23, 8'd232}: color_data = 12'ha00;
			{9'd23, 8'd233}: color_data = 12'ha00;
			{9'd23, 8'd234}: color_data = 12'h400;
			{9'd23, 8'd235}: color_data = 12'h510;
			{9'd23, 8'd236}: color_data = 12'hf40;
			{9'd23, 8'd237}: color_data = 12'hd10;
			{9'd23, 8'd238}: color_data = 12'h800;
			{9'd23, 8'd239}: color_data = 12'h100;
			{9'd24, 8'd16}: color_data = 12'h010;
			{9'd24, 8'd17}: color_data = 12'h780;
			{9'd24, 8'd18}: color_data = 12'hac0;
			{9'd24, 8'd19}: color_data = 12'hdea;
			{9'd24, 8'd20}: color_data = 12'hfff;
			{9'd24, 8'd21}: color_data = 12'hcd7;
			{9'd24, 8'd22}: color_data = 12'h9b0;
			{9'd24, 8'd23}: color_data = 12'h9b0;
			{9'd24, 8'd24}: color_data = 12'h9b0;
			{9'd24, 8'd25}: color_data = 12'h8a0;
			{9'd24, 8'd26}: color_data = 12'h450;
			{9'd24, 8'd27}: color_data = 12'h020;
			{9'd24, 8'd28}: color_data = 12'h140;
			{9'd24, 8'd29}: color_data = 12'h240;
			{9'd24, 8'd30}: color_data = 12'h660;
			{9'd24, 8'd31}: color_data = 12'h660;
			{9'd24, 8'd32}: color_data = 12'h110;
			{9'd24, 8'd68}: color_data = 12'h047;
			{9'd24, 8'd69}: color_data = 12'h6df;
			{9'd24, 8'd70}: color_data = 12'hfff;
			{9'd24, 8'd71}: color_data = 12'hfff;
			{9'd24, 8'd72}: color_data = 12'h9aa;
			{9'd24, 8'd73}: color_data = 12'h011;
			{9'd24, 8'd75}: color_data = 12'h012;
			{9'd24, 8'd76}: color_data = 12'h08c;
			{9'd24, 8'd77}: color_data = 12'h034;
			{9'd24, 8'd128}: color_data = 12'h047;
			{9'd24, 8'd129}: color_data = 12'h6df;
			{9'd24, 8'd130}: color_data = 12'hfff;
			{9'd24, 8'd131}: color_data = 12'hfff;
			{9'd24, 8'd132}: color_data = 12'h9aa;
			{9'd24, 8'd133}: color_data = 12'h111;
			{9'd24, 8'd135}: color_data = 12'h012;
			{9'd24, 8'd136}: color_data = 12'h08c;
			{9'd24, 8'd137}: color_data = 12'h034;
			{9'd24, 8'd170}: color_data = 12'h000;
			{9'd24, 8'd171}: color_data = 12'h068;
			{9'd24, 8'd172}: color_data = 12'h7ef;
			{9'd24, 8'd173}: color_data = 12'hfff;
			{9'd24, 8'd174}: color_data = 12'hfff;
			{9'd24, 8'd175}: color_data = 12'h899;
			{9'd24, 8'd176}: color_data = 12'h001;
			{9'd24, 8'd178}: color_data = 12'h024;
			{9'd24, 8'd179}: color_data = 12'h08c;
			{9'd24, 8'd180}: color_data = 12'h023;
			{9'd24, 8'd222}: color_data = 12'h200;
			{9'd24, 8'd223}: color_data = 12'h800;
			{9'd24, 8'd224}: color_data = 12'ha00;
			{9'd24, 8'd225}: color_data = 12'h800;
			{9'd24, 8'd226}: color_data = 12'h200;
			{9'd24, 8'd227}: color_data = 12'h920;
			{9'd24, 8'd228}: color_data = 12'hd30;
			{9'd24, 8'd229}: color_data = 12'h910;
			{9'd24, 8'd230}: color_data = 12'h200;
			{9'd24, 8'd231}: color_data = 12'h400;
			{9'd24, 8'd232}: color_data = 12'h900;
			{9'd24, 8'd233}: color_data = 12'ha00;
			{9'd24, 8'd234}: color_data = 12'h400;
			{9'd24, 8'd235}: color_data = 12'h310;
			{9'd24, 8'd236}: color_data = 12'hc30;
			{9'd24, 8'd237}: color_data = 12'hc20;
			{9'd24, 8'd238}: color_data = 12'h600;
			{9'd24, 8'd239}: color_data = 12'h000;
			{9'd25, 8'd16}: color_data = 12'h010;
			{9'd25, 8'd17}: color_data = 12'h780;
			{9'd25, 8'd18}: color_data = 12'hac0;
			{9'd25, 8'd19}: color_data = 12'hdea;
			{9'd25, 8'd20}: color_data = 12'hfff;
			{9'd25, 8'd21}: color_data = 12'hcd7;
			{9'd25, 8'd22}: color_data = 12'h9b0;
			{9'd25, 8'd23}: color_data = 12'h9b0;
			{9'd25, 8'd24}: color_data = 12'h9b0;
			{9'd25, 8'd25}: color_data = 12'h8a0;
			{9'd25, 8'd26}: color_data = 12'h450;
			{9'd25, 8'd27}: color_data = 12'h020;
			{9'd25, 8'd28}: color_data = 12'h140;
			{9'd25, 8'd29}: color_data = 12'h240;
			{9'd25, 8'd30}: color_data = 12'h660;
			{9'd25, 8'd31}: color_data = 12'h660;
			{9'd25, 8'd32}: color_data = 12'h110;
			{9'd25, 8'd68}: color_data = 12'h047;
			{9'd25, 8'd69}: color_data = 12'h6df;
			{9'd25, 8'd70}: color_data = 12'hfff;
			{9'd25, 8'd71}: color_data = 12'hcbb;
			{9'd25, 8'd72}: color_data = 12'h323;
			{9'd25, 8'd73}: color_data = 12'h002;
			{9'd25, 8'd74}: color_data = 12'h000;
			{9'd25, 8'd75}: color_data = 12'h012;
			{9'd25, 8'd76}: color_data = 12'h08c;
			{9'd25, 8'd77}: color_data = 12'h034;
			{9'd25, 8'd128}: color_data = 12'h047;
			{9'd25, 8'd129}: color_data = 12'h6df;
			{9'd25, 8'd130}: color_data = 12'hfff;
			{9'd25, 8'd131}: color_data = 12'hcbb;
			{9'd25, 8'd132}: color_data = 12'h323;
			{9'd25, 8'd133}: color_data = 12'h002;
			{9'd25, 8'd134}: color_data = 12'h000;
			{9'd25, 8'd135}: color_data = 12'h012;
			{9'd25, 8'd136}: color_data = 12'h08c;
			{9'd25, 8'd137}: color_data = 12'h034;
			{9'd25, 8'd170}: color_data = 12'h000;
			{9'd25, 8'd171}: color_data = 12'h068;
			{9'd25, 8'd172}: color_data = 12'h8ef;
			{9'd25, 8'd173}: color_data = 12'hfff;
			{9'd25, 8'd174}: color_data = 12'haaa;
			{9'd25, 8'd175}: color_data = 12'h213;
			{9'd25, 8'd176}: color_data = 12'h002;
			{9'd25, 8'd178}: color_data = 12'h023;
			{9'd25, 8'd179}: color_data = 12'h08c;
			{9'd25, 8'd180}: color_data = 12'h023;
			{9'd25, 8'd222}: color_data = 12'h200;
			{9'd25, 8'd223}: color_data = 12'h900;
			{9'd25, 8'd224}: color_data = 12'ha00;
			{9'd25, 8'd225}: color_data = 12'h800;
			{9'd25, 8'd226}: color_data = 12'h100;
			{9'd25, 8'd227}: color_data = 12'h100;
			{9'd25, 8'd228}: color_data = 12'h310;
			{9'd25, 8'd229}: color_data = 12'h200;
			{9'd25, 8'd230}: color_data = 12'h000;
			{9'd25, 8'd231}: color_data = 12'h500;
			{9'd25, 8'd232}: color_data = 12'ha00;
			{9'd25, 8'd233}: color_data = 12'ha00;
			{9'd25, 8'd234}: color_data = 12'h500;
			{9'd25, 8'd235}: color_data = 12'h000;
			{9'd25, 8'd236}: color_data = 12'h200;
			{9'd25, 8'd237}: color_data = 12'h300;
			{9'd25, 8'd238}: color_data = 12'h100;
			{9'd25, 8'd239}: color_data = 12'h000;
			{9'd26, 8'd16}: color_data = 12'h010;
			{9'd26, 8'd17}: color_data = 12'h780;
			{9'd26, 8'd18}: color_data = 12'hac0;
			{9'd26, 8'd19}: color_data = 12'hdea;
			{9'd26, 8'd20}: color_data = 12'hfff;
			{9'd26, 8'd21}: color_data = 12'hcd7;
			{9'd26, 8'd22}: color_data = 12'h9b0;
			{9'd26, 8'd23}: color_data = 12'h9b0;
			{9'd26, 8'd24}: color_data = 12'h9b0;
			{9'd26, 8'd25}: color_data = 12'h8a0;
			{9'd26, 8'd26}: color_data = 12'h450;
			{9'd26, 8'd27}: color_data = 12'h020;
			{9'd26, 8'd28}: color_data = 12'h140;
			{9'd26, 8'd29}: color_data = 12'h240;
			{9'd26, 8'd30}: color_data = 12'h660;
			{9'd26, 8'd31}: color_data = 12'h660;
			{9'd26, 8'd32}: color_data = 12'h110;
			{9'd26, 8'd68}: color_data = 12'h047;
			{9'd26, 8'd69}: color_data = 12'h6ef;
			{9'd26, 8'd70}: color_data = 12'hdcc;
			{9'd26, 8'd71}: color_data = 12'h434;
			{9'd26, 8'd72}: color_data = 12'h003;
			{9'd26, 8'd73}: color_data = 12'h005;
			{9'd26, 8'd74}: color_data = 12'h002;
			{9'd26, 8'd75}: color_data = 12'h012;
			{9'd26, 8'd76}: color_data = 12'h08c;
			{9'd26, 8'd77}: color_data = 12'h034;
			{9'd26, 8'd128}: color_data = 12'h047;
			{9'd26, 8'd129}: color_data = 12'h6ef;
			{9'd26, 8'd130}: color_data = 12'hddc;
			{9'd26, 8'd131}: color_data = 12'h434;
			{9'd26, 8'd132}: color_data = 12'h003;
			{9'd26, 8'd133}: color_data = 12'h005;
			{9'd26, 8'd134}: color_data = 12'h002;
			{9'd26, 8'd135}: color_data = 12'h012;
			{9'd26, 8'd136}: color_data = 12'h08c;
			{9'd26, 8'd137}: color_data = 12'h034;
			{9'd26, 8'd170}: color_data = 12'h000;
			{9'd26, 8'd171}: color_data = 12'h068;
			{9'd26, 8'd172}: color_data = 12'h8ff;
			{9'd26, 8'd173}: color_data = 12'hcbb;
			{9'd26, 8'd174}: color_data = 12'h323;
			{9'd26, 8'd175}: color_data = 12'h003;
			{9'd26, 8'd176}: color_data = 12'h005;
			{9'd26, 8'd177}: color_data = 12'h002;
			{9'd26, 8'd178}: color_data = 12'h023;
			{9'd26, 8'd179}: color_data = 12'h09c;
			{9'd26, 8'd180}: color_data = 12'h023;
			{9'd26, 8'd222}: color_data = 12'h300;
			{9'd26, 8'd223}: color_data = 12'hc20;
			{9'd26, 8'd224}: color_data = 12'ha00;
			{9'd26, 8'd225}: color_data = 12'h800;
			{9'd26, 8'd226}: color_data = 12'h100;
			{9'd26, 8'd227}: color_data = 12'h300;
			{9'd26, 8'd228}: color_data = 12'h500;
			{9'd26, 8'd229}: color_data = 12'h500;
			{9'd26, 8'd230}: color_data = 12'h100;
			{9'd26, 8'd231}: color_data = 12'h710;
			{9'd26, 8'd232}: color_data = 12'hc10;
			{9'd26, 8'd233}: color_data = 12'h900;
			{9'd26, 8'd234}: color_data = 12'h500;
			{9'd26, 8'd235}: color_data = 12'h100;
			{9'd26, 8'd236}: color_data = 12'h500;
			{9'd26, 8'd237}: color_data = 12'h500;
			{9'd26, 8'd238}: color_data = 12'h400;
			{9'd26, 8'd239}: color_data = 12'h000;
			{9'd27, 8'd16}: color_data = 12'h010;
			{9'd27, 8'd17}: color_data = 12'h780;
			{9'd27, 8'd18}: color_data = 12'hac0;
			{9'd27, 8'd19}: color_data = 12'hdea;
			{9'd27, 8'd20}: color_data = 12'hfff;
			{9'd27, 8'd21}: color_data = 12'hcd7;
			{9'd27, 8'd22}: color_data = 12'h9b0;
			{9'd27, 8'd23}: color_data = 12'h9b0;
			{9'd27, 8'd24}: color_data = 12'h9b0;
			{9'd27, 8'd25}: color_data = 12'h8a0;
			{9'd27, 8'd26}: color_data = 12'h450;
			{9'd27, 8'd27}: color_data = 12'h020;
			{9'd27, 8'd28}: color_data = 12'h140;
			{9'd27, 8'd29}: color_data = 12'h240;
			{9'd27, 8'd30}: color_data = 12'h660;
			{9'd27, 8'd31}: color_data = 12'h660;
			{9'd27, 8'd32}: color_data = 12'h110;
			{9'd27, 8'd68}: color_data = 12'h057;
			{9'd27, 8'd69}: color_data = 12'h3bd;
			{9'd27, 8'd70}: color_data = 12'h555;
			{9'd27, 8'd71}: color_data = 12'h002;
			{9'd27, 8'd72}: color_data = 12'h005;
			{9'd27, 8'd73}: color_data = 12'h005;
			{9'd27, 8'd74}: color_data = 12'h004;
			{9'd27, 8'd75}: color_data = 12'h025;
			{9'd27, 8'd76}: color_data = 12'h09c;
			{9'd27, 8'd77}: color_data = 12'h034;
			{9'd27, 8'd128}: color_data = 12'h057;
			{9'd27, 8'd129}: color_data = 12'h3bd;
			{9'd27, 8'd130}: color_data = 12'h555;
			{9'd27, 8'd131}: color_data = 12'h002;
			{9'd27, 8'd132}: color_data = 12'h005;
			{9'd27, 8'd133}: color_data = 12'h005;
			{9'd27, 8'd134}: color_data = 12'h004;
			{9'd27, 8'd135}: color_data = 12'h024;
			{9'd27, 8'd136}: color_data = 12'h09c;
			{9'd27, 8'd137}: color_data = 12'h034;
			{9'd27, 8'd170}: color_data = 12'h000;
			{9'd27, 8'd171}: color_data = 12'h079;
			{9'd27, 8'd172}: color_data = 12'h4bd;
			{9'd27, 8'd173}: color_data = 12'h444;
			{9'd27, 8'd174}: color_data = 12'h002;
			{9'd27, 8'd175}: color_data = 12'h005;
			{9'd27, 8'd176}: color_data = 12'h005;
			{9'd27, 8'd177}: color_data = 12'h004;
			{9'd27, 8'd178}: color_data = 12'h036;
			{9'd27, 8'd179}: color_data = 12'h09c;
			{9'd27, 8'd180}: color_data = 12'h023;
			{9'd27, 8'd222}: color_data = 12'h410;
			{9'd27, 8'd223}: color_data = 12'hd30;
			{9'd27, 8'd224}: color_data = 12'hb00;
			{9'd27, 8'd225}: color_data = 12'h700;
			{9'd27, 8'd226}: color_data = 12'h200;
			{9'd27, 8'd227}: color_data = 12'h700;
			{9'd27, 8'd228}: color_data = 12'hb00;
			{9'd27, 8'd229}: color_data = 12'ha00;
			{9'd27, 8'd230}: color_data = 12'h300;
			{9'd27, 8'd231}: color_data = 12'h820;
			{9'd27, 8'd232}: color_data = 12'hd20;
			{9'd27, 8'd233}: color_data = 12'h900;
			{9'd27, 8'd234}: color_data = 12'h500;
			{9'd27, 8'd235}: color_data = 12'h300;
			{9'd27, 8'd236}: color_data = 12'h900;
			{9'd27, 8'd237}: color_data = 12'hb00;
			{9'd27, 8'd238}: color_data = 12'h800;
			{9'd27, 8'd239}: color_data = 12'h100;
			{9'd28, 8'd16}: color_data = 12'h010;
			{9'd28, 8'd17}: color_data = 12'h780;
			{9'd28, 8'd18}: color_data = 12'hac0;
			{9'd28, 8'd19}: color_data = 12'hdea;
			{9'd28, 8'd20}: color_data = 12'hfff;
			{9'd28, 8'd21}: color_data = 12'hcd7;
			{9'd28, 8'd22}: color_data = 12'h9b0;
			{9'd28, 8'd23}: color_data = 12'h9b0;
			{9'd28, 8'd24}: color_data = 12'h9b0;
			{9'd28, 8'd25}: color_data = 12'h8a0;
			{9'd28, 8'd26}: color_data = 12'h450;
			{9'd28, 8'd27}: color_data = 12'h020;
			{9'd28, 8'd28}: color_data = 12'h140;
			{9'd28, 8'd29}: color_data = 12'h240;
			{9'd28, 8'd30}: color_data = 12'h660;
			{9'd28, 8'd31}: color_data = 12'h660;
			{9'd28, 8'd32}: color_data = 12'h110;
			{9'd28, 8'd68}: color_data = 12'h036;
			{9'd28, 8'd69}: color_data = 12'h047;
			{9'd28, 8'd70}: color_data = 12'h001;
			{9'd28, 8'd71}: color_data = 12'h004;
			{9'd28, 8'd72}: color_data = 12'h004;
			{9'd28, 8'd73}: color_data = 12'h004;
			{9'd28, 8'd74}: color_data = 12'h004;
			{9'd28, 8'd75}: color_data = 12'h015;
			{9'd28, 8'd76}: color_data = 12'h059;
			{9'd28, 8'd77}: color_data = 12'h023;
			{9'd28, 8'd128}: color_data = 12'h035;
			{9'd28, 8'd129}: color_data = 12'h047;
			{9'd28, 8'd130}: color_data = 12'h001;
			{9'd28, 8'd131}: color_data = 12'h004;
			{9'd28, 8'd132}: color_data = 12'h004;
			{9'd28, 8'd133}: color_data = 12'h004;
			{9'd28, 8'd134}: color_data = 12'h004;
			{9'd28, 8'd135}: color_data = 12'h015;
			{9'd28, 8'd136}: color_data = 12'h059;
			{9'd28, 8'd137}: color_data = 12'h023;
			{9'd28, 8'd170}: color_data = 12'h000;
			{9'd28, 8'd171}: color_data = 12'h047;
			{9'd28, 8'd172}: color_data = 12'h036;
			{9'd28, 8'd173}: color_data = 12'h001;
			{9'd28, 8'd174}: color_data = 12'h004;
			{9'd28, 8'd175}: color_data = 12'h004;
			{9'd28, 8'd176}: color_data = 12'h004;
			{9'd28, 8'd177}: color_data = 12'h004;
			{9'd28, 8'd178}: color_data = 12'h016;
			{9'd28, 8'd179}: color_data = 12'h059;
			{9'd28, 8'd180}: color_data = 12'h012;
			{9'd28, 8'd222}: color_data = 12'h410;
			{9'd28, 8'd223}: color_data = 12'he40;
			{9'd28, 8'd224}: color_data = 12'hd20;
			{9'd28, 8'd225}: color_data = 12'h800;
			{9'd28, 8'd226}: color_data = 12'h200;
			{9'd28, 8'd227}: color_data = 12'h700;
			{9'd28, 8'd228}: color_data = 12'hb00;
			{9'd28, 8'd229}: color_data = 12'h900;
			{9'd28, 8'd230}: color_data = 12'h300;
			{9'd28, 8'd231}: color_data = 12'h820;
			{9'd28, 8'd232}: color_data = 12'hf30;
			{9'd28, 8'd233}: color_data = 12'hc00;
			{9'd28, 8'd234}: color_data = 12'h500;
			{9'd28, 8'd235}: color_data = 12'h300;
			{9'd28, 8'd236}: color_data = 12'h900;
			{9'd28, 8'd237}: color_data = 12'hb00;
			{9'd28, 8'd238}: color_data = 12'h800;
			{9'd28, 8'd239}: color_data = 12'h100;
			{9'd29, 8'd16}: color_data = 12'h010;
			{9'd29, 8'd17}: color_data = 12'h780;
			{9'd29, 8'd18}: color_data = 12'hac0;
			{9'd29, 8'd19}: color_data = 12'hdea;
			{9'd29, 8'd20}: color_data = 12'hfff;
			{9'd29, 8'd21}: color_data = 12'hcd7;
			{9'd29, 8'd22}: color_data = 12'h9b0;
			{9'd29, 8'd23}: color_data = 12'h9b0;
			{9'd29, 8'd24}: color_data = 12'h9b0;
			{9'd29, 8'd25}: color_data = 12'h8a0;
			{9'd29, 8'd26}: color_data = 12'h450;
			{9'd29, 8'd27}: color_data = 12'h020;
			{9'd29, 8'd28}: color_data = 12'h140;
			{9'd29, 8'd29}: color_data = 12'h240;
			{9'd29, 8'd30}: color_data = 12'h660;
			{9'd29, 8'd31}: color_data = 12'h660;
			{9'd29, 8'd32}: color_data = 12'h110;
			{9'd29, 8'd68}: color_data = 12'h013;
			{9'd29, 8'd69}: color_data = 12'h027;
			{9'd29, 8'd70}: color_data = 12'h016;
			{9'd29, 8'd71}: color_data = 12'h027;
			{9'd29, 8'd72}: color_data = 12'h027;
			{9'd29, 8'd73}: color_data = 12'h027;
			{9'd29, 8'd74}: color_data = 12'h027;
			{9'd29, 8'd75}: color_data = 12'h028;
			{9'd29, 8'd76}: color_data = 12'h027;
			{9'd29, 8'd77}: color_data = 12'h001;
			{9'd29, 8'd128}: color_data = 12'h013;
			{9'd29, 8'd129}: color_data = 12'h027;
			{9'd29, 8'd130}: color_data = 12'h016;
			{9'd29, 8'd131}: color_data = 12'h027;
			{9'd29, 8'd132}: color_data = 12'h027;
			{9'd29, 8'd133}: color_data = 12'h026;
			{9'd29, 8'd134}: color_data = 12'h027;
			{9'd29, 8'd135}: color_data = 12'h028;
			{9'd29, 8'd136}: color_data = 12'h027;
			{9'd29, 8'd137}: color_data = 12'h001;
			{9'd29, 8'd170}: color_data = 12'h000;
			{9'd29, 8'd171}: color_data = 12'h014;
			{9'd29, 8'd172}: color_data = 12'h027;
			{9'd29, 8'd173}: color_data = 12'h016;
			{9'd29, 8'd174}: color_data = 12'h027;
			{9'd29, 8'd175}: color_data = 12'h027;
			{9'd29, 8'd176}: color_data = 12'h027;
			{9'd29, 8'd177}: color_data = 12'h027;
			{9'd29, 8'd178}: color_data = 12'h028;
			{9'd29, 8'd179}: color_data = 12'h026;
			{9'd29, 8'd180}: color_data = 12'h001;
			{9'd29, 8'd222}: color_data = 12'h310;
			{9'd29, 8'd223}: color_data = 12'he40;
			{9'd29, 8'd224}: color_data = 12'hc10;
			{9'd29, 8'd225}: color_data = 12'h800;
			{9'd29, 8'd226}: color_data = 12'h100;
			{9'd29, 8'd227}: color_data = 12'h700;
			{9'd29, 8'd228}: color_data = 12'ha00;
			{9'd29, 8'd229}: color_data = 12'ha00;
			{9'd29, 8'd230}: color_data = 12'h300;
			{9'd29, 8'd231}: color_data = 12'h720;
			{9'd29, 8'd232}: color_data = 12'he30;
			{9'd29, 8'd233}: color_data = 12'ha00;
			{9'd29, 8'd234}: color_data = 12'h600;
			{9'd29, 8'd235}: color_data = 12'h200;
			{9'd29, 8'd236}: color_data = 12'h900;
			{9'd29, 8'd237}: color_data = 12'ha00;
			{9'd29, 8'd238}: color_data = 12'h800;
			{9'd29, 8'd239}: color_data = 12'h100;
			{9'd30, 8'd16}: color_data = 12'h010;
			{9'd30, 8'd17}: color_data = 12'h780;
			{9'd30, 8'd18}: color_data = 12'hac0;
			{9'd30, 8'd19}: color_data = 12'hdea;
			{9'd30, 8'd20}: color_data = 12'hfff;
			{9'd30, 8'd21}: color_data = 12'hcd7;
			{9'd30, 8'd22}: color_data = 12'h9b0;
			{9'd30, 8'd23}: color_data = 12'h9b0;
			{9'd30, 8'd24}: color_data = 12'h9c0;
			{9'd30, 8'd25}: color_data = 12'h8a0;
			{9'd30, 8'd26}: color_data = 12'h450;
			{9'd30, 8'd27}: color_data = 12'h020;
			{9'd30, 8'd28}: color_data = 12'h140;
			{9'd30, 8'd29}: color_data = 12'h240;
			{9'd30, 8'd30}: color_data = 12'h660;
			{9'd30, 8'd31}: color_data = 12'h660;
			{9'd30, 8'd32}: color_data = 12'h110;
			{9'd30, 8'd68}: color_data = 12'h036;
			{9'd30, 8'd69}: color_data = 12'h09e;
			{9'd30, 8'd70}: color_data = 12'h09e;
			{9'd30, 8'd71}: color_data = 12'h09e;
			{9'd30, 8'd72}: color_data = 12'h09e;
			{9'd30, 8'd73}: color_data = 12'h09e;
			{9'd30, 8'd74}: color_data = 12'h09e;
			{9'd30, 8'd75}: color_data = 12'h09e;
			{9'd30, 8'd76}: color_data = 12'h08c;
			{9'd30, 8'd77}: color_data = 12'h023;
			{9'd30, 8'd128}: color_data = 12'h035;
			{9'd30, 8'd129}: color_data = 12'h09e;
			{9'd30, 8'd130}: color_data = 12'h09e;
			{9'd30, 8'd131}: color_data = 12'h09e;
			{9'd30, 8'd132}: color_data = 12'h09e;
			{9'd30, 8'd133}: color_data = 12'h09e;
			{9'd30, 8'd134}: color_data = 12'h09e;
			{9'd30, 8'd135}: color_data = 12'h09e;
			{9'd30, 8'd136}: color_data = 12'h08c;
			{9'd30, 8'd137}: color_data = 12'h023;
			{9'd30, 8'd170}: color_data = 12'h000;
			{9'd30, 8'd171}: color_data = 12'h057;
			{9'd30, 8'd172}: color_data = 12'h0ae;
			{9'd30, 8'd173}: color_data = 12'h09e;
			{9'd30, 8'd174}: color_data = 12'h09e;
			{9'd30, 8'd175}: color_data = 12'h09e;
			{9'd30, 8'd176}: color_data = 12'h09e;
			{9'd30, 8'd177}: color_data = 12'h09e;
			{9'd30, 8'd178}: color_data = 12'h09e;
			{9'd30, 8'd179}: color_data = 12'h07b;
			{9'd30, 8'd180}: color_data = 12'h012;
			{9'd30, 8'd222}: color_data = 12'h310;
			{9'd30, 8'd223}: color_data = 12'he30;
			{9'd30, 8'd224}: color_data = 12'hb10;
			{9'd30, 8'd225}: color_data = 12'h900;
			{9'd30, 8'd226}: color_data = 12'h100;
			{9'd30, 8'd227}: color_data = 12'h600;
			{9'd30, 8'd228}: color_data = 12'ha00;
			{9'd30, 8'd229}: color_data = 12'ha00;
			{9'd30, 8'd230}: color_data = 12'h300;
			{9'd30, 8'd231}: color_data = 12'h720;
			{9'd30, 8'd232}: color_data = 12'he30;
			{9'd30, 8'd233}: color_data = 12'ha00;
			{9'd30, 8'd234}: color_data = 12'h700;
			{9'd30, 8'd235}: color_data = 12'h100;
			{9'd30, 8'd236}: color_data = 12'h800;
			{9'd30, 8'd237}: color_data = 12'ha00;
			{9'd30, 8'd238}: color_data = 12'h800;
			{9'd30, 8'd239}: color_data = 12'h000;
			{9'd31, 8'd16}: color_data = 12'h010;
			{9'd31, 8'd17}: color_data = 12'h780;
			{9'd31, 8'd18}: color_data = 12'hac0;
			{9'd31, 8'd19}: color_data = 12'hdea;
			{9'd31, 8'd20}: color_data = 12'hfff;
			{9'd31, 8'd21}: color_data = 12'hcd7;
			{9'd31, 8'd22}: color_data = 12'h9b0;
			{9'd31, 8'd23}: color_data = 12'h9b0;
			{9'd31, 8'd24}: color_data = 12'h9c0;
			{9'd31, 8'd25}: color_data = 12'h9a0;
			{9'd31, 8'd26}: color_data = 12'h450;
			{9'd31, 8'd27}: color_data = 12'h020;
			{9'd31, 8'd28}: color_data = 12'h140;
			{9'd31, 8'd29}: color_data = 12'h240;
			{9'd31, 8'd30}: color_data = 12'h660;
			{9'd31, 8'd31}: color_data = 12'h660;
			{9'd31, 8'd32}: color_data = 12'h110;
			{9'd31, 8'd68}: color_data = 12'h057;
			{9'd31, 8'd69}: color_data = 12'h4ef;
			{9'd31, 8'd70}: color_data = 12'h7ef;
			{9'd31, 8'd71}: color_data = 12'h0cf;
			{9'd31, 8'd72}: color_data = 12'h0cf;
			{9'd31, 8'd73}: color_data = 12'h0df;
			{9'd31, 8'd74}: color_data = 12'h0bd;
			{9'd31, 8'd75}: color_data = 12'h068;
			{9'd31, 8'd76}: color_data = 12'h09c;
			{9'd31, 8'd77}: color_data = 12'h034;
			{9'd31, 8'd128}: color_data = 12'h057;
			{9'd31, 8'd129}: color_data = 12'h4ef;
			{9'd31, 8'd130}: color_data = 12'h7ef;
			{9'd31, 8'd131}: color_data = 12'h0cf;
			{9'd31, 8'd132}: color_data = 12'h0cf;
			{9'd31, 8'd133}: color_data = 12'h0df;
			{9'd31, 8'd134}: color_data = 12'h0bd;
			{9'd31, 8'd135}: color_data = 12'h068;
			{9'd31, 8'd136}: color_data = 12'h09c;
			{9'd31, 8'd137}: color_data = 12'h034;
			{9'd31, 8'd170}: color_data = 12'h000;
			{9'd31, 8'd171}: color_data = 12'h069;
			{9'd31, 8'd172}: color_data = 12'h6ef;
			{9'd31, 8'd173}: color_data = 12'h6ef;
			{9'd31, 8'd174}: color_data = 12'h0cf;
			{9'd31, 8'd175}: color_data = 12'h0cf;
			{9'd31, 8'd176}: color_data = 12'h0df;
			{9'd31, 8'd177}: color_data = 12'h0ac;
			{9'd31, 8'd178}: color_data = 12'h079;
			{9'd31, 8'd179}: color_data = 12'h09c;
			{9'd31, 8'd180}: color_data = 12'h023;
			{9'd31, 8'd222}: color_data = 12'h300;
			{9'd31, 8'd223}: color_data = 12'he40;
			{9'd31, 8'd224}: color_data = 12'he30;
			{9'd31, 8'd225}: color_data = 12'h900;
			{9'd31, 8'd226}: color_data = 12'h100;
			{9'd31, 8'd227}: color_data = 12'h600;
			{9'd31, 8'd228}: color_data = 12'ha00;
			{9'd31, 8'd229}: color_data = 12'h900;
			{9'd31, 8'd230}: color_data = 12'h300;
			{9'd31, 8'd231}: color_data = 12'h620;
			{9'd31, 8'd232}: color_data = 12'hf40;
			{9'd31, 8'd233}: color_data = 12'hd20;
			{9'd31, 8'd234}: color_data = 12'h600;
			{9'd31, 8'd235}: color_data = 12'h100;
			{9'd31, 8'd236}: color_data = 12'h800;
			{9'd31, 8'd237}: color_data = 12'ha00;
			{9'd31, 8'd238}: color_data = 12'h800;
			{9'd31, 8'd239}: color_data = 12'h000;
			{9'd32, 8'd16}: color_data = 12'h000;
			{9'd32, 8'd17}: color_data = 12'h660;
			{9'd32, 8'd18}: color_data = 12'h890;
			{9'd32, 8'd19}: color_data = 12'hdda;
			{9'd32, 8'd20}: color_data = 12'hfff;
			{9'd32, 8'd21}: color_data = 12'hbc7;
			{9'd32, 8'd22}: color_data = 12'h780;
			{9'd32, 8'd23}: color_data = 12'h890;
			{9'd32, 8'd24}: color_data = 12'h890;
			{9'd32, 8'd25}: color_data = 12'h880;
			{9'd32, 8'd26}: color_data = 12'h450;
			{9'd32, 8'd27}: color_data = 12'h020;
			{9'd32, 8'd28}: color_data = 12'h140;
			{9'd32, 8'd29}: color_data = 12'h250;
			{9'd32, 8'd30}: color_data = 12'h660;
			{9'd32, 8'd31}: color_data = 12'h660;
			{9'd32, 8'd32}: color_data = 12'h110;
			{9'd32, 8'd68}: color_data = 12'h047;
			{9'd32, 8'd69}: color_data = 12'h6df;
			{9'd32, 8'd70}: color_data = 12'heff;
			{9'd32, 8'd71}: color_data = 12'h6df;
			{9'd32, 8'd72}: color_data = 12'h0bf;
			{9'd32, 8'd73}: color_data = 12'h0bf;
			{9'd32, 8'd74}: color_data = 12'h056;
			{9'd32, 8'd75}: color_data = 12'h012;
			{9'd32, 8'd76}: color_data = 12'h08b;
			{9'd32, 8'd77}: color_data = 12'h034;
			{9'd32, 8'd128}: color_data = 12'h047;
			{9'd32, 8'd129}: color_data = 12'h6df;
			{9'd32, 8'd130}: color_data = 12'heff;
			{9'd32, 8'd131}: color_data = 12'h6df;
			{9'd32, 8'd132}: color_data = 12'h0bf;
			{9'd32, 8'd133}: color_data = 12'h0bf;
			{9'd32, 8'd134}: color_data = 12'h056;
			{9'd32, 8'd135}: color_data = 12'h012;
			{9'd32, 8'd136}: color_data = 12'h08b;
			{9'd32, 8'd137}: color_data = 12'h034;
			{9'd32, 8'd170}: color_data = 12'h000;
			{9'd32, 8'd171}: color_data = 12'h068;
			{9'd32, 8'd172}: color_data = 12'h8ef;
			{9'd32, 8'd173}: color_data = 12'hdff;
			{9'd32, 8'd174}: color_data = 12'h4cf;
			{9'd32, 8'd175}: color_data = 12'h0cf;
			{9'd32, 8'd176}: color_data = 12'h0ae;
			{9'd32, 8'd177}: color_data = 12'h035;
			{9'd32, 8'd178}: color_data = 12'h023;
			{9'd32, 8'd179}: color_data = 12'h08c;
			{9'd32, 8'd180}: color_data = 12'h023;
			{9'd32, 8'd222}: color_data = 12'h000;
			{9'd32, 8'd223}: color_data = 12'h410;
			{9'd32, 8'd224}: color_data = 12'h410;
			{9'd32, 8'd225}: color_data = 12'h200;
			{9'd32, 8'd226}: color_data = 12'h000;
			{9'd32, 8'd227}: color_data = 12'h600;
			{9'd32, 8'd228}: color_data = 12'h900;
			{9'd32, 8'd229}: color_data = 12'h900;
			{9'd32, 8'd230}: color_data = 12'h400;
			{9'd32, 8'd231}: color_data = 12'h100;
			{9'd32, 8'd232}: color_data = 12'h410;
			{9'd32, 8'd233}: color_data = 12'h410;
			{9'd32, 8'd234}: color_data = 12'h100;
			{9'd32, 8'd235}: color_data = 12'h100;
			{9'd32, 8'd236}: color_data = 12'h800;
			{9'd32, 8'd237}: color_data = 12'ha00;
			{9'd32, 8'd238}: color_data = 12'h800;
			{9'd32, 8'd239}: color_data = 12'h000;
			{9'd33, 8'd16}: color_data = 12'h000;
			{9'd33, 8'd17}: color_data = 12'h230;
			{9'd33, 8'd18}: color_data = 12'h340;
			{9'd33, 8'd19}: color_data = 12'h786;
			{9'd33, 8'd20}: color_data = 12'habb;
			{9'd33, 8'd21}: color_data = 12'h674;
			{9'd33, 8'd22}: color_data = 12'h330;
			{9'd33, 8'd23}: color_data = 12'h340;
			{9'd33, 8'd24}: color_data = 12'h340;
			{9'd33, 8'd25}: color_data = 12'h340;
			{9'd33, 8'd26}: color_data = 12'h230;
			{9'd33, 8'd27}: color_data = 12'h020;
			{9'd33, 8'd28}: color_data = 12'h030;
			{9'd33, 8'd29}: color_data = 12'h130;
			{9'd33, 8'd30}: color_data = 12'h440;
			{9'd33, 8'd31}: color_data = 12'h340;
			{9'd33, 8'd32}: color_data = 12'h010;
			{9'd33, 8'd68}: color_data = 12'h047;
			{9'd33, 8'd69}: color_data = 12'h6df;
			{9'd33, 8'd70}: color_data = 12'hfff;
			{9'd33, 8'd71}: color_data = 12'hdff;
			{9'd33, 8'd72}: color_data = 12'h5df;
			{9'd33, 8'd73}: color_data = 12'h068;
			{9'd33, 8'd74}: color_data = 12'h000;
			{9'd33, 8'd75}: color_data = 12'h012;
			{9'd33, 8'd76}: color_data = 12'h08c;
			{9'd33, 8'd77}: color_data = 12'h034;
			{9'd33, 8'd128}: color_data = 12'h047;
			{9'd33, 8'd129}: color_data = 12'h6df;
			{9'd33, 8'd130}: color_data = 12'hfff;
			{9'd33, 8'd131}: color_data = 12'hdff;
			{9'd33, 8'd132}: color_data = 12'h5df;
			{9'd33, 8'd133}: color_data = 12'h068;
			{9'd33, 8'd134}: color_data = 12'h000;
			{9'd33, 8'd135}: color_data = 12'h012;
			{9'd33, 8'd136}: color_data = 12'h08c;
			{9'd33, 8'd137}: color_data = 12'h034;
			{9'd33, 8'd170}: color_data = 12'h000;
			{9'd33, 8'd171}: color_data = 12'h068;
			{9'd33, 8'd172}: color_data = 12'h8ef;
			{9'd33, 8'd173}: color_data = 12'hfff;
			{9'd33, 8'd174}: color_data = 12'hcff;
			{9'd33, 8'd175}: color_data = 12'h4ce;
			{9'd33, 8'd176}: color_data = 12'h057;
			{9'd33, 8'd177}: color_data = 12'h000;
			{9'd33, 8'd178}: color_data = 12'h023;
			{9'd33, 8'd179}: color_data = 12'h08c;
			{9'd33, 8'd180}: color_data = 12'h023;
			{9'd33, 8'd222}: color_data = 12'h000;
			{9'd33, 8'd223}: color_data = 12'h300;
			{9'd33, 8'd224}: color_data = 12'h300;
			{9'd33, 8'd225}: color_data = 12'h300;
			{9'd33, 8'd226}: color_data = 12'h100;
			{9'd33, 8'd227}: color_data = 12'h910;
			{9'd33, 8'd228}: color_data = 12'hb00;
			{9'd33, 8'd229}: color_data = 12'h900;
			{9'd33, 8'd230}: color_data = 12'h400;
			{9'd33, 8'd231}: color_data = 12'h100;
			{9'd33, 8'd232}: color_data = 12'h300;
			{9'd33, 8'd233}: color_data = 12'h400;
			{9'd33, 8'd234}: color_data = 12'h200;
			{9'd33, 8'd235}: color_data = 12'h200;
			{9'd33, 8'd236}: color_data = 12'hb10;
			{9'd33, 8'd237}: color_data = 12'ha00;
			{9'd33, 8'd238}: color_data = 12'h800;
			{9'd33, 8'd239}: color_data = 12'h000;
			{9'd34, 8'd15}: color_data = 12'h000;
			{9'd34, 8'd16}: color_data = 12'h110;
			{9'd34, 8'd17}: color_data = 12'h130;
			{9'd34, 8'd18}: color_data = 12'h242;
			{9'd34, 8'd19}: color_data = 12'h343;
			{9'd34, 8'd20}: color_data = 12'h242;
			{9'd34, 8'd21}: color_data = 12'h130;
			{9'd34, 8'd22}: color_data = 12'h130;
			{9'd34, 8'd23}: color_data = 12'h130;
			{9'd34, 8'd24}: color_data = 12'h130;
			{9'd34, 8'd25}: color_data = 12'h130;
			{9'd34, 8'd26}: color_data = 12'h130;
			{9'd34, 8'd27}: color_data = 12'h020;
			{9'd34, 8'd28}: color_data = 12'h020;
			{9'd34, 8'd29}: color_data = 12'h020;
			{9'd34, 8'd30}: color_data = 12'h020;
			{9'd34, 8'd31}: color_data = 12'h120;
			{9'd34, 8'd32}: color_data = 12'h110;
			{9'd34, 8'd33}: color_data = 12'h000;
			{9'd34, 8'd68}: color_data = 12'h047;
			{9'd34, 8'd69}: color_data = 12'h6df;
			{9'd34, 8'd70}: color_data = 12'hfff;
			{9'd34, 8'd71}: color_data = 12'hfff;
			{9'd34, 8'd72}: color_data = 12'h9aa;
			{9'd34, 8'd73}: color_data = 12'h011;
			{9'd34, 8'd75}: color_data = 12'h012;
			{9'd34, 8'd76}: color_data = 12'h08c;
			{9'd34, 8'd77}: color_data = 12'h034;
			{9'd34, 8'd128}: color_data = 12'h047;
			{9'd34, 8'd129}: color_data = 12'h6df;
			{9'd34, 8'd130}: color_data = 12'hfff;
			{9'd34, 8'd131}: color_data = 12'hfff;
			{9'd34, 8'd132}: color_data = 12'h9aa;
			{9'd34, 8'd133}: color_data = 12'h111;
			{9'd34, 8'd135}: color_data = 12'h012;
			{9'd34, 8'd136}: color_data = 12'h08c;
			{9'd34, 8'd137}: color_data = 12'h034;
			{9'd34, 8'd170}: color_data = 12'h000;
			{9'd34, 8'd171}: color_data = 12'h068;
			{9'd34, 8'd172}: color_data = 12'h7ef;
			{9'd34, 8'd173}: color_data = 12'hfff;
			{9'd34, 8'd174}: color_data = 12'hfff;
			{9'd34, 8'd175}: color_data = 12'h899;
			{9'd34, 8'd176}: color_data = 12'h001;
			{9'd34, 8'd178}: color_data = 12'h024;
			{9'd34, 8'd179}: color_data = 12'h08c;
			{9'd34, 8'd180}: color_data = 12'h023;
			{9'd34, 8'd222}: color_data = 12'h200;
			{9'd34, 8'd223}: color_data = 12'h900;
			{9'd34, 8'd224}: color_data = 12'ha00;
			{9'd34, 8'd225}: color_data = 12'h900;
			{9'd34, 8'd226}: color_data = 12'h200;
			{9'd34, 8'd227}: color_data = 12'hb30;
			{9'd34, 8'd228}: color_data = 12'hc10;
			{9'd34, 8'd229}: color_data = 12'h900;
			{9'd34, 8'd230}: color_data = 12'h300;
			{9'd34, 8'd231}: color_data = 12'h300;
			{9'd34, 8'd232}: color_data = 12'ha00;
			{9'd34, 8'd233}: color_data = 12'ha00;
			{9'd34, 8'd234}: color_data = 12'h600;
			{9'd34, 8'd235}: color_data = 12'h310;
			{9'd34, 8'd236}: color_data = 12'he30;
			{9'd34, 8'd237}: color_data = 12'ha00;
			{9'd34, 8'd238}: color_data = 12'h700;
			{9'd34, 8'd239}: color_data = 12'h000;
			{9'd35, 8'd15}: color_data = 12'h010;
			{9'd35, 8'd16}: color_data = 12'h670;
			{9'd35, 8'd17}: color_data = 12'h8a0;
			{9'd35, 8'd18}: color_data = 12'hbc9;
			{9'd35, 8'd19}: color_data = 12'hcdd;
			{9'd35, 8'd20}: color_data = 12'h9a4;
			{9'd35, 8'd21}: color_data = 12'h790;
			{9'd35, 8'd22}: color_data = 12'h790;
			{9'd35, 8'd23}: color_data = 12'h790;
			{9'd35, 8'd24}: color_data = 12'h790;
			{9'd35, 8'd25}: color_data = 12'h7a0;
			{9'd35, 8'd26}: color_data = 12'h780;
			{9'd35, 8'd27}: color_data = 12'h440;
			{9'd35, 8'd28}: color_data = 12'h020;
			{9'd35, 8'd29}: color_data = 12'h130;
			{9'd35, 8'd30}: color_data = 12'h140;
			{9'd35, 8'd31}: color_data = 12'h450;
			{9'd35, 8'd32}: color_data = 12'h550;
			{9'd35, 8'd33}: color_data = 12'h110;
			{9'd35, 8'd68}: color_data = 12'h047;
			{9'd35, 8'd69}: color_data = 12'h6df;
			{9'd35, 8'd70}: color_data = 12'hfff;
			{9'd35, 8'd71}: color_data = 12'hcbb;
			{9'd35, 8'd72}: color_data = 12'h323;
			{9'd35, 8'd73}: color_data = 12'h002;
			{9'd35, 8'd74}: color_data = 12'h000;
			{9'd35, 8'd75}: color_data = 12'h012;
			{9'd35, 8'd76}: color_data = 12'h08c;
			{9'd35, 8'd77}: color_data = 12'h034;
			{9'd35, 8'd128}: color_data = 12'h047;
			{9'd35, 8'd129}: color_data = 12'h6df;
			{9'd35, 8'd130}: color_data = 12'hfff;
			{9'd35, 8'd131}: color_data = 12'hcbb;
			{9'd35, 8'd132}: color_data = 12'h323;
			{9'd35, 8'd133}: color_data = 12'h002;
			{9'd35, 8'd134}: color_data = 12'h000;
			{9'd35, 8'd135}: color_data = 12'h012;
			{9'd35, 8'd136}: color_data = 12'h08c;
			{9'd35, 8'd137}: color_data = 12'h034;
			{9'd35, 8'd170}: color_data = 12'h000;
			{9'd35, 8'd171}: color_data = 12'h068;
			{9'd35, 8'd172}: color_data = 12'h8ef;
			{9'd35, 8'd173}: color_data = 12'hfff;
			{9'd35, 8'd174}: color_data = 12'haaa;
			{9'd35, 8'd175}: color_data = 12'h213;
			{9'd35, 8'd176}: color_data = 12'h002;
			{9'd35, 8'd177}: color_data = 12'h000;
			{9'd35, 8'd178}: color_data = 12'h023;
			{9'd35, 8'd179}: color_data = 12'h08c;
			{9'd35, 8'd180}: color_data = 12'h023;
			{9'd35, 8'd222}: color_data = 12'h200;
			{9'd35, 8'd223}: color_data = 12'h900;
			{9'd35, 8'd224}: color_data = 12'ha00;
			{9'd35, 8'd225}: color_data = 12'h800;
			{9'd35, 8'd226}: color_data = 12'h100;
			{9'd35, 8'd227}: color_data = 12'hb30;
			{9'd35, 8'd228}: color_data = 12'hd20;
			{9'd35, 8'd229}: color_data = 12'ha00;
			{9'd35, 8'd230}: color_data = 12'h400;
			{9'd35, 8'd231}: color_data = 12'h300;
			{9'd35, 8'd232}: color_data = 12'ha00;
			{9'd35, 8'd233}: color_data = 12'ha00;
			{9'd35, 8'd234}: color_data = 12'h600;
			{9'd35, 8'd235}: color_data = 12'h310;
			{9'd35, 8'd236}: color_data = 12'he40;
			{9'd35, 8'd237}: color_data = 12'hc10;
			{9'd35, 8'd238}: color_data = 12'h800;
			{9'd35, 8'd239}: color_data = 12'h000;
			{9'd36, 8'd15}: color_data = 12'h110;
			{9'd36, 8'd16}: color_data = 12'h890;
			{9'd36, 8'd17}: color_data = 12'had1;
			{9'd36, 8'd18}: color_data = 12'hefb;
			{9'd36, 8'd19}: color_data = 12'hfff;
			{9'd36, 8'd20}: color_data = 12'hcd6;
			{9'd36, 8'd21}: color_data = 12'h9b0;
			{9'd36, 8'd22}: color_data = 12'hac0;
			{9'd36, 8'd23}: color_data = 12'hac0;
			{9'd36, 8'd24}: color_data = 12'hac0;
			{9'd36, 8'd25}: color_data = 12'hac0;
			{9'd36, 8'd26}: color_data = 12'h9b0;
			{9'd36, 8'd27}: color_data = 12'h550;
			{9'd36, 8'd28}: color_data = 12'h020;
			{9'd36, 8'd29}: color_data = 12'h140;
			{9'd36, 8'd30}: color_data = 12'h240;
			{9'd36, 8'd31}: color_data = 12'h660;
			{9'd36, 8'd32}: color_data = 12'h760;
			{9'd36, 8'd33}: color_data = 12'h120;
			{9'd36, 8'd68}: color_data = 12'h047;
			{9'd36, 8'd69}: color_data = 12'h6ef;
			{9'd36, 8'd70}: color_data = 12'hddc;
			{9'd36, 8'd71}: color_data = 12'h434;
			{9'd36, 8'd72}: color_data = 12'h003;
			{9'd36, 8'd73}: color_data = 12'h005;
			{9'd36, 8'd74}: color_data = 12'h002;
			{9'd36, 8'd75}: color_data = 12'h012;
			{9'd36, 8'd76}: color_data = 12'h08c;
			{9'd36, 8'd77}: color_data = 12'h034;
			{9'd36, 8'd128}: color_data = 12'h047;
			{9'd36, 8'd129}: color_data = 12'h6ef;
			{9'd36, 8'd130}: color_data = 12'hddc;
			{9'd36, 8'd131}: color_data = 12'h434;
			{9'd36, 8'd132}: color_data = 12'h003;
			{9'd36, 8'd133}: color_data = 12'h005;
			{9'd36, 8'd134}: color_data = 12'h002;
			{9'd36, 8'd135}: color_data = 12'h012;
			{9'd36, 8'd136}: color_data = 12'h08c;
			{9'd36, 8'd137}: color_data = 12'h034;
			{9'd36, 8'd170}: color_data = 12'h000;
			{9'd36, 8'd171}: color_data = 12'h068;
			{9'd36, 8'd172}: color_data = 12'h8ff;
			{9'd36, 8'd173}: color_data = 12'hcbb;
			{9'd36, 8'd174}: color_data = 12'h323;
			{9'd36, 8'd175}: color_data = 12'h003;
			{9'd36, 8'd176}: color_data = 12'h005;
			{9'd36, 8'd177}: color_data = 12'h002;
			{9'd36, 8'd178}: color_data = 12'h023;
			{9'd36, 8'd179}: color_data = 12'h09c;
			{9'd36, 8'd180}: color_data = 12'h023;
			{9'd36, 8'd222}: color_data = 12'h200;
			{9'd36, 8'd223}: color_data = 12'h800;
			{9'd36, 8'd224}: color_data = 12'ha00;
			{9'd36, 8'd225}: color_data = 12'h800;
			{9'd36, 8'd226}: color_data = 12'h100;
			{9'd36, 8'd227}: color_data = 12'ha30;
			{9'd36, 8'd228}: color_data = 12'hf40;
			{9'd36, 8'd229}: color_data = 12'hb10;
			{9'd36, 8'd230}: color_data = 12'h300;
			{9'd36, 8'd231}: color_data = 12'h300;
			{9'd36, 8'd232}: color_data = 12'h900;
			{9'd36, 8'd233}: color_data = 12'ha00;
			{9'd36, 8'd234}: color_data = 12'h600;
			{9'd36, 8'd235}: color_data = 12'h200;
			{9'd36, 8'd236}: color_data = 12'hd40;
			{9'd36, 8'd237}: color_data = 12'he30;
			{9'd36, 8'd238}: color_data = 12'h800;
			{9'd36, 8'd239}: color_data = 12'h000;
			{9'd37, 8'd15}: color_data = 12'h110;
			{9'd37, 8'd16}: color_data = 12'h790;
			{9'd37, 8'd17}: color_data = 12'h9c0;
			{9'd37, 8'd18}: color_data = 12'heeb;
			{9'd37, 8'd19}: color_data = 12'hfff;
			{9'd37, 8'd20}: color_data = 12'hbd6;
			{9'd37, 8'd21}: color_data = 12'h8b0;
			{9'd37, 8'd22}: color_data = 12'h9b0;
			{9'd37, 8'd23}: color_data = 12'h9b0;
			{9'd37, 8'd24}: color_data = 12'h9b0;
			{9'd37, 8'd25}: color_data = 12'h9b0;
			{9'd37, 8'd26}: color_data = 12'h9a0;
			{9'd37, 8'd27}: color_data = 12'h550;
			{9'd37, 8'd28}: color_data = 12'h020;
			{9'd37, 8'd29}: color_data = 12'h130;
			{9'd37, 8'd30}: color_data = 12'h240;
			{9'd37, 8'd31}: color_data = 12'h660;
			{9'd37, 8'd32}: color_data = 12'h660;
			{9'd37, 8'd33}: color_data = 12'h110;
			{9'd37, 8'd68}: color_data = 12'h057;
			{9'd37, 8'd69}: color_data = 12'h3bd;
			{9'd37, 8'd70}: color_data = 12'h555;
			{9'd37, 8'd71}: color_data = 12'h002;
			{9'd37, 8'd72}: color_data = 12'h005;
			{9'd37, 8'd73}: color_data = 12'h005;
			{9'd37, 8'd74}: color_data = 12'h004;
			{9'd37, 8'd75}: color_data = 12'h025;
			{9'd37, 8'd76}: color_data = 12'h09c;
			{9'd37, 8'd77}: color_data = 12'h034;
			{9'd37, 8'd128}: color_data = 12'h057;
			{9'd37, 8'd129}: color_data = 12'h3bd;
			{9'd37, 8'd130}: color_data = 12'h555;
			{9'd37, 8'd131}: color_data = 12'h002;
			{9'd37, 8'd132}: color_data = 12'h005;
			{9'd37, 8'd133}: color_data = 12'h005;
			{9'd37, 8'd134}: color_data = 12'h004;
			{9'd37, 8'd135}: color_data = 12'h025;
			{9'd37, 8'd136}: color_data = 12'h09c;
			{9'd37, 8'd137}: color_data = 12'h034;
			{9'd37, 8'd170}: color_data = 12'h000;
			{9'd37, 8'd171}: color_data = 12'h079;
			{9'd37, 8'd172}: color_data = 12'h4bd;
			{9'd37, 8'd173}: color_data = 12'h444;
			{9'd37, 8'd174}: color_data = 12'h002;
			{9'd37, 8'd175}: color_data = 12'h005;
			{9'd37, 8'd176}: color_data = 12'h005;
			{9'd37, 8'd177}: color_data = 12'h004;
			{9'd37, 8'd178}: color_data = 12'h036;
			{9'd37, 8'd179}: color_data = 12'h09c;
			{9'd37, 8'd180}: color_data = 12'h023;
			{9'd37, 8'd222}: color_data = 12'h100;
			{9'd37, 8'd223}: color_data = 12'h800;
			{9'd37, 8'd224}: color_data = 12'ha00;
			{9'd37, 8'd225}: color_data = 12'h900;
			{9'd37, 8'd226}: color_data = 12'h100;
			{9'd37, 8'd227}: color_data = 12'h200;
			{9'd37, 8'd228}: color_data = 12'h410;
			{9'd37, 8'd229}: color_data = 12'h200;
			{9'd37, 8'd230}: color_data = 12'h000;
			{9'd37, 8'd231}: color_data = 12'h300;
			{9'd37, 8'd232}: color_data = 12'h900;
			{9'd37, 8'd233}: color_data = 12'ha00;
			{9'd37, 8'd234}: color_data = 12'h700;
			{9'd37, 8'd235}: color_data = 12'h000;
			{9'd37, 8'd236}: color_data = 12'h310;
			{9'd37, 8'd237}: color_data = 12'h410;
			{9'd37, 8'd238}: color_data = 12'h200;
			{9'd38, 8'd15}: color_data = 12'h110;
			{9'd38, 8'd16}: color_data = 12'h8a0;
			{9'd38, 8'd17}: color_data = 12'hce5;
			{9'd38, 8'd18}: color_data = 12'hffd;
			{9'd38, 8'd19}: color_data = 12'hfff;
			{9'd38, 8'd20}: color_data = 12'heea;
			{9'd38, 8'd21}: color_data = 12'hbc2;
			{9'd38, 8'd22}: color_data = 12'h9c0;
			{9'd38, 8'd23}: color_data = 12'hac0;
			{9'd38, 8'd24}: color_data = 12'hac0;
			{9'd38, 8'd25}: color_data = 12'hac0;
			{9'd38, 8'd26}: color_data = 12'h9b0;
			{9'd38, 8'd27}: color_data = 12'h550;
			{9'd38, 8'd28}: color_data = 12'h020;
			{9'd38, 8'd29}: color_data = 12'h140;
			{9'd38, 8'd30}: color_data = 12'h250;
			{9'd38, 8'd31}: color_data = 12'h660;
			{9'd38, 8'd32}: color_data = 12'h760;
			{9'd38, 8'd33}: color_data = 12'h110;
			{9'd38, 8'd68}: color_data = 12'h036;
			{9'd38, 8'd69}: color_data = 12'h047;
			{9'd38, 8'd70}: color_data = 12'h001;
			{9'd38, 8'd71}: color_data = 12'h004;
			{9'd38, 8'd72}: color_data = 12'h004;
			{9'd38, 8'd73}: color_data = 12'h004;
			{9'd38, 8'd74}: color_data = 12'h004;
			{9'd38, 8'd75}: color_data = 12'h015;
			{9'd38, 8'd76}: color_data = 12'h059;
			{9'd38, 8'd77}: color_data = 12'h023;
			{9'd38, 8'd128}: color_data = 12'h036;
			{9'd38, 8'd129}: color_data = 12'h058;
			{9'd38, 8'd130}: color_data = 12'h002;
			{9'd38, 8'd131}: color_data = 12'h005;
			{9'd38, 8'd132}: color_data = 12'h005;
			{9'd38, 8'd133}: color_data = 12'h005;
			{9'd38, 8'd134}: color_data = 12'h005;
			{9'd38, 8'd135}: color_data = 12'h017;
			{9'd38, 8'd136}: color_data = 12'h05a;
			{9'd38, 8'd137}: color_data = 12'h023;
			{9'd38, 8'd170}: color_data = 12'h000;
			{9'd38, 8'd171}: color_data = 12'h047;
			{9'd38, 8'd172}: color_data = 12'h036;
			{9'd38, 8'd173}: color_data = 12'h001;
			{9'd38, 8'd174}: color_data = 12'h004;
			{9'd38, 8'd175}: color_data = 12'h004;
			{9'd38, 8'd176}: color_data = 12'h004;
			{9'd38, 8'd177}: color_data = 12'h004;
			{9'd38, 8'd178}: color_data = 12'h016;
			{9'd38, 8'd179}: color_data = 12'h059;
			{9'd38, 8'd180}: color_data = 12'h012;
			{9'd38, 8'd222}: color_data = 12'h200;
			{9'd38, 8'd223}: color_data = 12'hc20;
			{9'd38, 8'd224}: color_data = 12'ha00;
			{9'd38, 8'd225}: color_data = 12'h800;
			{9'd38, 8'd226}: color_data = 12'h100;
			{9'd38, 8'd227}: color_data = 12'h200;
			{9'd38, 8'd228}: color_data = 12'h400;
			{9'd38, 8'd229}: color_data = 12'h400;
			{9'd38, 8'd230}: color_data = 12'h100;
			{9'd38, 8'd231}: color_data = 12'h510;
			{9'd38, 8'd232}: color_data = 12'hc10;
			{9'd38, 8'd233}: color_data = 12'ha00;
			{9'd38, 8'd234}: color_data = 12'h700;
			{9'd38, 8'd235}: color_data = 12'h000;
			{9'd38, 8'd236}: color_data = 12'h300;
			{9'd38, 8'd237}: color_data = 12'h400;
			{9'd38, 8'd238}: color_data = 12'h300;
			{9'd38, 8'd239}: color_data = 12'h000;
			{9'd39, 8'd15}: color_data = 12'h010;
			{9'd39, 8'd16}: color_data = 12'h681;
			{9'd39, 8'd17}: color_data = 12'hcd9;
			{9'd39, 8'd18}: color_data = 12'hddd;
			{9'd39, 8'd19}: color_data = 12'hddd;
			{9'd39, 8'd20}: color_data = 12'hddd;
			{9'd39, 8'd21}: color_data = 12'hab5;
			{9'd39, 8'd22}: color_data = 12'h790;
			{9'd39, 8'd23}: color_data = 12'h790;
			{9'd39, 8'd24}: color_data = 12'h790;
			{9'd39, 8'd25}: color_data = 12'h890;
			{9'd39, 8'd26}: color_data = 12'h780;
			{9'd39, 8'd27}: color_data = 12'h440;
			{9'd39, 8'd28}: color_data = 12'h020;
			{9'd39, 8'd29}: color_data = 12'h130;
			{9'd39, 8'd30}: color_data = 12'h230;
			{9'd39, 8'd31}: color_data = 12'h550;
			{9'd39, 8'd32}: color_data = 12'h550;
			{9'd39, 8'd33}: color_data = 12'h110;
			{9'd39, 8'd68}: color_data = 12'h013;
			{9'd39, 8'd69}: color_data = 12'h027;
			{9'd39, 8'd70}: color_data = 12'h016;
			{9'd39, 8'd71}: color_data = 12'h027;
			{9'd39, 8'd72}: color_data = 12'h027;
			{9'd39, 8'd73}: color_data = 12'h017;
			{9'd39, 8'd74}: color_data = 12'h027;
			{9'd39, 8'd75}: color_data = 12'h028;
			{9'd39, 8'd76}: color_data = 12'h027;
			{9'd39, 8'd77}: color_data = 12'h001;
			{9'd39, 8'd128}: color_data = 12'h002;
			{9'd39, 8'd129}: color_data = 12'h004;
			{9'd39, 8'd130}: color_data = 12'h004;
			{9'd39, 8'd131}: color_data = 12'h004;
			{9'd39, 8'd132}: color_data = 12'h004;
			{9'd39, 8'd133}: color_data = 12'h004;
			{9'd39, 8'd134}: color_data = 12'h004;
			{9'd39, 8'd135}: color_data = 12'h004;
			{9'd39, 8'd136}: color_data = 12'h004;
			{9'd39, 8'd137}: color_data = 12'h001;
			{9'd39, 8'd170}: color_data = 12'h000;
			{9'd39, 8'd171}: color_data = 12'h014;
			{9'd39, 8'd172}: color_data = 12'h027;
			{9'd39, 8'd173}: color_data = 12'h016;
			{9'd39, 8'd174}: color_data = 12'h027;
			{9'd39, 8'd175}: color_data = 12'h027;
			{9'd39, 8'd176}: color_data = 12'h016;
			{9'd39, 8'd177}: color_data = 12'h027;
			{9'd39, 8'd178}: color_data = 12'h028;
			{9'd39, 8'd179}: color_data = 12'h026;
			{9'd39, 8'd180}: color_data = 12'h001;
			{9'd39, 8'd222}: color_data = 12'h310;
			{9'd39, 8'd223}: color_data = 12'he30;
			{9'd39, 8'd224}: color_data = 12'ha00;
			{9'd39, 8'd225}: color_data = 12'h800;
			{9'd39, 8'd226}: color_data = 12'h100;
			{9'd39, 8'd227}: color_data = 12'h600;
			{9'd39, 8'd228}: color_data = 12'ha00;
			{9'd39, 8'd229}: color_data = 12'ha00;
			{9'd39, 8'd230}: color_data = 12'h300;
			{9'd39, 8'd231}: color_data = 12'h720;
			{9'd39, 8'd232}: color_data = 12'he30;
			{9'd39, 8'd233}: color_data = 12'h900;
			{9'd39, 8'd234}: color_data = 12'h600;
			{9'd39, 8'd235}: color_data = 12'h100;
			{9'd39, 8'd236}: color_data = 12'h900;
			{9'd39, 8'd237}: color_data = 12'ha00;
			{9'd39, 8'd238}: color_data = 12'h800;
			{9'd39, 8'd239}: color_data = 12'h000;
			{9'd40, 8'd15}: color_data = 12'h000;
			{9'd40, 8'd16}: color_data = 12'h110;
			{9'd40, 8'd17}: color_data = 12'h222;
			{9'd40, 8'd18}: color_data = 12'h323;
			{9'd40, 8'd19}: color_data = 12'h222;
			{9'd40, 8'd20}: color_data = 12'h333;
			{9'd40, 8'd21}: color_data = 12'h221;
			{9'd40, 8'd22}: color_data = 12'h120;
			{9'd40, 8'd23}: color_data = 12'h120;
			{9'd40, 8'd24}: color_data = 12'h120;
			{9'd40, 8'd25}: color_data = 12'h120;
			{9'd40, 8'd26}: color_data = 12'h110;
			{9'd40, 8'd27}: color_data = 12'h000;
			{9'd40, 8'd28}: color_data = 12'h000;
			{9'd40, 8'd29}: color_data = 12'h000;
			{9'd40, 8'd30}: color_data = 12'h000;
			{9'd40, 8'd31}: color_data = 12'h110;
			{9'd40, 8'd32}: color_data = 12'h110;
			{9'd40, 8'd33}: color_data = 12'h000;
			{9'd40, 8'd68}: color_data = 12'h035;
			{9'd40, 8'd69}: color_data = 12'h09e;
			{9'd40, 8'd70}: color_data = 12'h09e;
			{9'd40, 8'd71}: color_data = 12'h09e;
			{9'd40, 8'd72}: color_data = 12'h09e;
			{9'd40, 8'd73}: color_data = 12'h09e;
			{9'd40, 8'd74}: color_data = 12'h09e;
			{9'd40, 8'd75}: color_data = 12'h09e;
			{9'd40, 8'd76}: color_data = 12'h08c;
			{9'd40, 8'd77}: color_data = 12'h023;
			{9'd40, 8'd128}: color_data = 12'h000;
			{9'd40, 8'd129}: color_data = 12'h000;
			{9'd40, 8'd130}: color_data = 12'h001;
			{9'd40, 8'd131}: color_data = 12'h001;
			{9'd40, 8'd132}: color_data = 12'h000;
			{9'd40, 8'd133}: color_data = 12'h000;
			{9'd40, 8'd134}: color_data = 12'h000;
			{9'd40, 8'd135}: color_data = 12'h000;
			{9'd40, 8'd136}: color_data = 12'h000;
			{9'd40, 8'd137}: color_data = 12'h000;
			{9'd40, 8'd170}: color_data = 12'h000;
			{9'd40, 8'd171}: color_data = 12'h057;
			{9'd40, 8'd172}: color_data = 12'h0ae;
			{9'd40, 8'd173}: color_data = 12'h09e;
			{9'd40, 8'd174}: color_data = 12'h09e;
			{9'd40, 8'd175}: color_data = 12'h09e;
			{9'd40, 8'd176}: color_data = 12'h09e;
			{9'd40, 8'd177}: color_data = 12'h09e;
			{9'd40, 8'd178}: color_data = 12'h09e;
			{9'd40, 8'd179}: color_data = 12'h07b;
			{9'd40, 8'd180}: color_data = 12'h012;
			{9'd40, 8'd222}: color_data = 12'h310;
			{9'd40, 8'd223}: color_data = 12'he40;
			{9'd40, 8'd224}: color_data = 12'hc10;
			{9'd40, 8'd225}: color_data = 12'h900;
			{9'd40, 8'd226}: color_data = 12'h100;
			{9'd40, 8'd227}: color_data = 12'h600;
			{9'd40, 8'd228}: color_data = 12'ha00;
			{9'd40, 8'd229}: color_data = 12'ha00;
			{9'd40, 8'd230}: color_data = 12'h300;
			{9'd40, 8'd231}: color_data = 12'h720;
			{9'd40, 8'd232}: color_data = 12'hf30;
			{9'd40, 8'd233}: color_data = 12'hb00;
			{9'd40, 8'd234}: color_data = 12'h700;
			{9'd40, 8'd235}: color_data = 12'h100;
			{9'd40, 8'd236}: color_data = 12'h800;
			{9'd40, 8'd237}: color_data = 12'ha00;
			{9'd40, 8'd238}: color_data = 12'h800;
			{9'd40, 8'd239}: color_data = 12'h000;
			{9'd41, 8'd68}: color_data = 12'h057;
			{9'd41, 8'd69}: color_data = 12'h4ef;
			{9'd41, 8'd70}: color_data = 12'h7ef;
			{9'd41, 8'd71}: color_data = 12'h0cf;
			{9'd41, 8'd72}: color_data = 12'h0cf;
			{9'd41, 8'd73}: color_data = 12'h0df;
			{9'd41, 8'd74}: color_data = 12'h0bd;
			{9'd41, 8'd75}: color_data = 12'h068;
			{9'd41, 8'd76}: color_data = 12'h09c;
			{9'd41, 8'd77}: color_data = 12'h034;
			{9'd41, 8'd170}: color_data = 12'h000;
			{9'd41, 8'd171}: color_data = 12'h069;
			{9'd41, 8'd172}: color_data = 12'h6ef;
			{9'd41, 8'd173}: color_data = 12'h6ef;
			{9'd41, 8'd174}: color_data = 12'h0cf;
			{9'd41, 8'd175}: color_data = 12'h0cf;
			{9'd41, 8'd176}: color_data = 12'h0df;
			{9'd41, 8'd177}: color_data = 12'h0ad;
			{9'd41, 8'd178}: color_data = 12'h079;
			{9'd41, 8'd179}: color_data = 12'h09c;
			{9'd41, 8'd180}: color_data = 12'h023;
			{9'd41, 8'd222}: color_data = 12'h300;
			{9'd41, 8'd223}: color_data = 12'hd40;
			{9'd41, 8'd224}: color_data = 12'he30;
			{9'd41, 8'd225}: color_data = 12'h800;
			{9'd41, 8'd226}: color_data = 12'h100;
			{9'd41, 8'd227}: color_data = 12'h600;
			{9'd41, 8'd228}: color_data = 12'ha00;
			{9'd41, 8'd229}: color_data = 12'h900;
			{9'd41, 8'd230}: color_data = 12'h300;
			{9'd41, 8'd231}: color_data = 12'h610;
			{9'd41, 8'd232}: color_data = 12'hf40;
			{9'd41, 8'd233}: color_data = 12'hd20;
			{9'd41, 8'd234}: color_data = 12'h600;
			{9'd41, 8'd235}: color_data = 12'h100;
			{9'd41, 8'd236}: color_data = 12'h800;
			{9'd41, 8'd237}: color_data = 12'ha00;
			{9'd41, 8'd238}: color_data = 12'h800;
			{9'd41, 8'd239}: color_data = 12'h000;
			{9'd42, 8'd68}: color_data = 12'h047;
			{9'd42, 8'd69}: color_data = 12'h6df;
			{9'd42, 8'd70}: color_data = 12'heff;
			{9'd42, 8'd71}: color_data = 12'h6df;
			{9'd42, 8'd72}: color_data = 12'h0bf;
			{9'd42, 8'd73}: color_data = 12'h0be;
			{9'd42, 8'd74}: color_data = 12'h056;
			{9'd42, 8'd75}: color_data = 12'h012;
			{9'd42, 8'd76}: color_data = 12'h08b;
			{9'd42, 8'd77}: color_data = 12'h034;
			{9'd42, 8'd170}: color_data = 12'h000;
			{9'd42, 8'd171}: color_data = 12'h068;
			{9'd42, 8'd172}: color_data = 12'h8ef;
			{9'd42, 8'd173}: color_data = 12'hdff;
			{9'd42, 8'd174}: color_data = 12'h4cf;
			{9'd42, 8'd175}: color_data = 12'h0bf;
			{9'd42, 8'd176}: color_data = 12'h0ae;
			{9'd42, 8'd177}: color_data = 12'h035;
			{9'd42, 8'd178}: color_data = 12'h023;
			{9'd42, 8'd179}: color_data = 12'h08c;
			{9'd42, 8'd180}: color_data = 12'h023;
			{9'd42, 8'd222}: color_data = 12'h000;
			{9'd42, 8'd223}: color_data = 12'h310;
			{9'd42, 8'd224}: color_data = 12'h310;
			{9'd42, 8'd225}: color_data = 12'h100;
			{9'd42, 8'd226}: color_data = 12'h000;
			{9'd42, 8'd227}: color_data = 12'h600;
			{9'd42, 8'd228}: color_data = 12'ha00;
			{9'd42, 8'd229}: color_data = 12'h900;
			{9'd42, 8'd230}: color_data = 12'h400;
			{9'd42, 8'd231}: color_data = 12'h000;
			{9'd42, 8'd232}: color_data = 12'h310;
			{9'd42, 8'd233}: color_data = 12'h300;
			{9'd42, 8'd234}: color_data = 12'h000;
			{9'd42, 8'd235}: color_data = 12'h100;
			{9'd42, 8'd236}: color_data = 12'h800;
			{9'd42, 8'd237}: color_data = 12'ha00;
			{9'd42, 8'd238}: color_data = 12'h800;
			{9'd42, 8'd239}: color_data = 12'h000;
			{9'd43, 8'd68}: color_data = 12'h047;
			{9'd43, 8'd69}: color_data = 12'h6df;
			{9'd43, 8'd70}: color_data = 12'hfff;
			{9'd43, 8'd71}: color_data = 12'hdff;
			{9'd43, 8'd72}: color_data = 12'h5df;
			{9'd43, 8'd73}: color_data = 12'h068;
			{9'd43, 8'd74}: color_data = 12'h000;
			{9'd43, 8'd75}: color_data = 12'h012;
			{9'd43, 8'd76}: color_data = 12'h08c;
			{9'd43, 8'd77}: color_data = 12'h034;
			{9'd43, 8'd170}: color_data = 12'h000;
			{9'd43, 8'd171}: color_data = 12'h068;
			{9'd43, 8'd172}: color_data = 12'h8ef;
			{9'd43, 8'd173}: color_data = 12'hfff;
			{9'd43, 8'd174}: color_data = 12'hcff;
			{9'd43, 8'd175}: color_data = 12'h4ce;
			{9'd43, 8'd176}: color_data = 12'h057;
			{9'd43, 8'd177}: color_data = 12'h000;
			{9'd43, 8'd178}: color_data = 12'h023;
			{9'd43, 8'd179}: color_data = 12'h08c;
			{9'd43, 8'd180}: color_data = 12'h023;
			{9'd43, 8'd222}: color_data = 12'h100;
			{9'd43, 8'd223}: color_data = 12'h400;
			{9'd43, 8'd224}: color_data = 12'h500;
			{9'd43, 8'd225}: color_data = 12'h400;
			{9'd43, 8'd226}: color_data = 12'h100;
			{9'd43, 8'd227}: color_data = 12'h920;
			{9'd43, 8'd228}: color_data = 12'hb10;
			{9'd43, 8'd229}: color_data = 12'h900;
			{9'd43, 8'd230}: color_data = 12'h400;
			{9'd43, 8'd231}: color_data = 12'h100;
			{9'd43, 8'd232}: color_data = 12'h400;
			{9'd43, 8'd233}: color_data = 12'h500;
			{9'd43, 8'd234}: color_data = 12'h300;
			{9'd43, 8'd235}: color_data = 12'h200;
			{9'd43, 8'd236}: color_data = 12'hc20;
			{9'd43, 8'd237}: color_data = 12'ha00;
			{9'd43, 8'd238}: color_data = 12'h800;
			{9'd43, 8'd239}: color_data = 12'h000;
			{9'd44, 8'd68}: color_data = 12'h047;
			{9'd44, 8'd69}: color_data = 12'h6df;
			{9'd44, 8'd70}: color_data = 12'hfff;
			{9'd44, 8'd71}: color_data = 12'hfff;
			{9'd44, 8'd72}: color_data = 12'h9aa;
			{9'd44, 8'd73}: color_data = 12'h011;
			{9'd44, 8'd75}: color_data = 12'h012;
			{9'd44, 8'd76}: color_data = 12'h08c;
			{9'd44, 8'd77}: color_data = 12'h034;
			{9'd44, 8'd170}: color_data = 12'h000;
			{9'd44, 8'd171}: color_data = 12'h068;
			{9'd44, 8'd172}: color_data = 12'h7ef;
			{9'd44, 8'd173}: color_data = 12'hfff;
			{9'd44, 8'd174}: color_data = 12'hfff;
			{9'd44, 8'd175}: color_data = 12'h899;
			{9'd44, 8'd176}: color_data = 12'h001;
			{9'd44, 8'd178}: color_data = 12'h024;
			{9'd44, 8'd179}: color_data = 12'h08c;
			{9'd44, 8'd180}: color_data = 12'h023;
			{9'd44, 8'd222}: color_data = 12'h200;
			{9'd44, 8'd223}: color_data = 12'h900;
			{9'd44, 8'd224}: color_data = 12'ha00;
			{9'd44, 8'd225}: color_data = 12'h900;
			{9'd44, 8'd226}: color_data = 12'h200;
			{9'd44, 8'd227}: color_data = 12'hb30;
			{9'd44, 8'd228}: color_data = 12'hc10;
			{9'd44, 8'd229}: color_data = 12'h900;
			{9'd44, 8'd230}: color_data = 12'h300;
			{9'd44, 8'd231}: color_data = 12'h300;
			{9'd44, 8'd232}: color_data = 12'ha00;
			{9'd44, 8'd233}: color_data = 12'ha00;
			{9'd44, 8'd234}: color_data = 12'h600;
			{9'd44, 8'd235}: color_data = 12'h310;
			{9'd44, 8'd236}: color_data = 12'he30;
			{9'd44, 8'd237}: color_data = 12'ha00;
			{9'd44, 8'd238}: color_data = 12'h700;
			{9'd44, 8'd239}: color_data = 12'h000;
			{9'd45, 8'd68}: color_data = 12'h047;
			{9'd45, 8'd69}: color_data = 12'h6df;
			{9'd45, 8'd70}: color_data = 12'hfff;
			{9'd45, 8'd71}: color_data = 12'hcbb;
			{9'd45, 8'd72}: color_data = 12'h323;
			{9'd45, 8'd73}: color_data = 12'h002;
			{9'd45, 8'd74}: color_data = 12'h000;
			{9'd45, 8'd75}: color_data = 12'h012;
			{9'd45, 8'd76}: color_data = 12'h08c;
			{9'd45, 8'd77}: color_data = 12'h034;
			{9'd45, 8'd170}: color_data = 12'h000;
			{9'd45, 8'd171}: color_data = 12'h068;
			{9'd45, 8'd172}: color_data = 12'h8ef;
			{9'd45, 8'd173}: color_data = 12'hfff;
			{9'd45, 8'd174}: color_data = 12'haaa;
			{9'd45, 8'd175}: color_data = 12'h213;
			{9'd45, 8'd176}: color_data = 12'h002;
			{9'd45, 8'd178}: color_data = 12'h023;
			{9'd45, 8'd179}: color_data = 12'h08c;
			{9'd45, 8'd180}: color_data = 12'h023;
			{9'd45, 8'd222}: color_data = 12'h200;
			{9'd45, 8'd223}: color_data = 12'h900;
			{9'd45, 8'd224}: color_data = 12'ha00;
			{9'd45, 8'd225}: color_data = 12'h800;
			{9'd45, 8'd226}: color_data = 12'h100;
			{9'd45, 8'd227}: color_data = 12'hb30;
			{9'd45, 8'd228}: color_data = 12'he20;
			{9'd45, 8'd229}: color_data = 12'ha00;
			{9'd45, 8'd230}: color_data = 12'h400;
			{9'd45, 8'd231}: color_data = 12'h300;
			{9'd45, 8'd232}: color_data = 12'h900;
			{9'd45, 8'd233}: color_data = 12'ha00;
			{9'd45, 8'd234}: color_data = 12'h600;
			{9'd45, 8'd235}: color_data = 12'h310;
			{9'd45, 8'd236}: color_data = 12'he40;
			{9'd45, 8'd237}: color_data = 12'hc10;
			{9'd45, 8'd238}: color_data = 12'h800;
			{9'd45, 8'd239}: color_data = 12'h000;
			{9'd46, 8'd68}: color_data = 12'h047;
			{9'd46, 8'd69}: color_data = 12'h6ef;
			{9'd46, 8'd70}: color_data = 12'hdcc;
			{9'd46, 8'd71}: color_data = 12'h434;
			{9'd46, 8'd72}: color_data = 12'h003;
			{9'd46, 8'd73}: color_data = 12'h005;
			{9'd46, 8'd74}: color_data = 12'h002;
			{9'd46, 8'd75}: color_data = 12'h012;
			{9'd46, 8'd76}: color_data = 12'h08c;
			{9'd46, 8'd77}: color_data = 12'h034;
			{9'd46, 8'd170}: color_data = 12'h000;
			{9'd46, 8'd171}: color_data = 12'h068;
			{9'd46, 8'd172}: color_data = 12'h8ff;
			{9'd46, 8'd173}: color_data = 12'hcbb;
			{9'd46, 8'd174}: color_data = 12'h323;
			{9'd46, 8'd175}: color_data = 12'h003;
			{9'd46, 8'd176}: color_data = 12'h005;
			{9'd46, 8'd177}: color_data = 12'h002;
			{9'd46, 8'd178}: color_data = 12'h023;
			{9'd46, 8'd179}: color_data = 12'h09c;
			{9'd46, 8'd180}: color_data = 12'h023;
			{9'd46, 8'd222}: color_data = 12'h100;
			{9'd46, 8'd223}: color_data = 12'h800;
			{9'd46, 8'd224}: color_data = 12'ha00;
			{9'd46, 8'd225}: color_data = 12'h800;
			{9'd46, 8'd226}: color_data = 12'h100;
			{9'd46, 8'd227}: color_data = 12'h930;
			{9'd46, 8'd228}: color_data = 12'he40;
			{9'd46, 8'd229}: color_data = 12'hb10;
			{9'd46, 8'd230}: color_data = 12'h300;
			{9'd46, 8'd231}: color_data = 12'h300;
			{9'd46, 8'd232}: color_data = 12'h900;
			{9'd46, 8'd233}: color_data = 12'ha00;
			{9'd46, 8'd234}: color_data = 12'h600;
			{9'd46, 8'd235}: color_data = 12'h200;
			{9'd46, 8'd236}: color_data = 12'hc30;
			{9'd46, 8'd237}: color_data = 12'he30;
			{9'd46, 8'd238}: color_data = 12'h800;
			{9'd46, 8'd239}: color_data = 12'h000;
			{9'd47, 8'd68}: color_data = 12'h057;
			{9'd47, 8'd69}: color_data = 12'h3bd;
			{9'd47, 8'd70}: color_data = 12'h555;
			{9'd47, 8'd71}: color_data = 12'h002;
			{9'd47, 8'd72}: color_data = 12'h005;
			{9'd47, 8'd73}: color_data = 12'h005;
			{9'd47, 8'd74}: color_data = 12'h004;
			{9'd47, 8'd75}: color_data = 12'h025;
			{9'd47, 8'd76}: color_data = 12'h09c;
			{9'd47, 8'd77}: color_data = 12'h034;
			{9'd47, 8'd170}: color_data = 12'h000;
			{9'd47, 8'd171}: color_data = 12'h079;
			{9'd47, 8'd172}: color_data = 12'h4bd;
			{9'd47, 8'd173}: color_data = 12'h444;
			{9'd47, 8'd174}: color_data = 12'h002;
			{9'd47, 8'd175}: color_data = 12'h005;
			{9'd47, 8'd176}: color_data = 12'h005;
			{9'd47, 8'd177}: color_data = 12'h004;
			{9'd47, 8'd178}: color_data = 12'h036;
			{9'd47, 8'd179}: color_data = 12'h09c;
			{9'd47, 8'd180}: color_data = 12'h023;
			{9'd47, 8'd222}: color_data = 12'h200;
			{9'd47, 8'd223}: color_data = 12'h900;
			{9'd47, 8'd224}: color_data = 12'ha00;
			{9'd47, 8'd225}: color_data = 12'h900;
			{9'd47, 8'd226}: color_data = 12'h100;
			{9'd47, 8'd227}: color_data = 12'h100;
			{9'd47, 8'd228}: color_data = 12'h310;
			{9'd47, 8'd229}: color_data = 12'h200;
			{9'd47, 8'd230}: color_data = 12'h000;
			{9'd47, 8'd231}: color_data = 12'h400;
			{9'd47, 8'd232}: color_data = 12'h900;
			{9'd47, 8'd233}: color_data = 12'ha00;
			{9'd47, 8'd234}: color_data = 12'h700;
			{9'd47, 8'd235}: color_data = 12'h000;
			{9'd47, 8'd236}: color_data = 12'h200;
			{9'd47, 8'd237}: color_data = 12'h210;
			{9'd47, 8'd238}: color_data = 12'h100;
			{9'd48, 8'd68}: color_data = 12'h036;
			{9'd48, 8'd69}: color_data = 12'h047;
			{9'd48, 8'd70}: color_data = 12'h001;
			{9'd48, 8'd71}: color_data = 12'h004;
			{9'd48, 8'd72}: color_data = 12'h004;
			{9'd48, 8'd73}: color_data = 12'h004;
			{9'd48, 8'd74}: color_data = 12'h004;
			{9'd48, 8'd75}: color_data = 12'h015;
			{9'd48, 8'd76}: color_data = 12'h059;
			{9'd48, 8'd77}: color_data = 12'h023;
			{9'd48, 8'd170}: color_data = 12'h000;
			{9'd48, 8'd171}: color_data = 12'h047;
			{9'd48, 8'd172}: color_data = 12'h036;
			{9'd48, 8'd173}: color_data = 12'h001;
			{9'd48, 8'd174}: color_data = 12'h004;
			{9'd48, 8'd175}: color_data = 12'h004;
			{9'd48, 8'd176}: color_data = 12'h004;
			{9'd48, 8'd177}: color_data = 12'h004;
			{9'd48, 8'd178}: color_data = 12'h016;
			{9'd48, 8'd179}: color_data = 12'h059;
			{9'd48, 8'd180}: color_data = 12'h012;
			{9'd48, 8'd222}: color_data = 12'h300;
			{9'd48, 8'd223}: color_data = 12'hc20;
			{9'd48, 8'd224}: color_data = 12'ha00;
			{9'd48, 8'd225}: color_data = 12'h800;
			{9'd48, 8'd226}: color_data = 12'h100;
			{9'd48, 8'd227}: color_data = 12'h300;
			{9'd48, 8'd228}: color_data = 12'h500;
			{9'd48, 8'd229}: color_data = 12'h500;
			{9'd48, 8'd230}: color_data = 12'h100;
			{9'd48, 8'd231}: color_data = 12'h610;
			{9'd48, 8'd232}: color_data = 12'hc20;
			{9'd48, 8'd233}: color_data = 12'ha00;
			{9'd48, 8'd234}: color_data = 12'h600;
			{9'd48, 8'd235}: color_data = 12'h100;
			{9'd48, 8'd236}: color_data = 12'h400;
			{9'd48, 8'd237}: color_data = 12'h500;
			{9'd48, 8'd238}: color_data = 12'h400;
			{9'd48, 8'd239}: color_data = 12'h000;
			{9'd49, 8'd68}: color_data = 12'h013;
			{9'd49, 8'd69}: color_data = 12'h027;
			{9'd49, 8'd70}: color_data = 12'h016;
			{9'd49, 8'd71}: color_data = 12'h027;
			{9'd49, 8'd72}: color_data = 12'h027;
			{9'd49, 8'd73}: color_data = 12'h026;
			{9'd49, 8'd74}: color_data = 12'h027;
			{9'd49, 8'd75}: color_data = 12'h028;
			{9'd49, 8'd76}: color_data = 12'h027;
			{9'd49, 8'd77}: color_data = 12'h001;
			{9'd49, 8'd170}: color_data = 12'h000;
			{9'd49, 8'd171}: color_data = 12'h014;
			{9'd49, 8'd172}: color_data = 12'h027;
			{9'd49, 8'd173}: color_data = 12'h016;
			{9'd49, 8'd174}: color_data = 12'h027;
			{9'd49, 8'd175}: color_data = 12'h027;
			{9'd49, 8'd176}: color_data = 12'h026;
			{9'd49, 8'd177}: color_data = 12'h027;
			{9'd49, 8'd178}: color_data = 12'h028;
			{9'd49, 8'd179}: color_data = 12'h026;
			{9'd49, 8'd180}: color_data = 12'h001;
			{9'd49, 8'd222}: color_data = 12'h310;
			{9'd49, 8'd223}: color_data = 12'he30;
			{9'd49, 8'd224}: color_data = 12'ha00;
			{9'd49, 8'd225}: color_data = 12'h800;
			{9'd49, 8'd226}: color_data = 12'h100;
			{9'd49, 8'd227}: color_data = 12'h700;
			{9'd49, 8'd228}: color_data = 12'ha00;
			{9'd49, 8'd229}: color_data = 12'ha00;
			{9'd49, 8'd230}: color_data = 12'h300;
			{9'd49, 8'd231}: color_data = 12'h720;
			{9'd49, 8'd232}: color_data = 12'he30;
			{9'd49, 8'd233}: color_data = 12'h900;
			{9'd49, 8'd234}: color_data = 12'h600;
			{9'd49, 8'd235}: color_data = 12'h100;
			{9'd49, 8'd236}: color_data = 12'h900;
			{9'd49, 8'd237}: color_data = 12'ha00;
			{9'd49, 8'd238}: color_data = 12'h800;
			{9'd49, 8'd239}: color_data = 12'h000;
			{9'd50, 8'd68}: color_data = 12'h035;
			{9'd50, 8'd69}: color_data = 12'h09e;
			{9'd50, 8'd70}: color_data = 12'h09e;
			{9'd50, 8'd71}: color_data = 12'h09e;
			{9'd50, 8'd72}: color_data = 12'h09e;
			{9'd50, 8'd73}: color_data = 12'h09e;
			{9'd50, 8'd74}: color_data = 12'h09e;
			{9'd50, 8'd75}: color_data = 12'h09e;
			{9'd50, 8'd76}: color_data = 12'h08c;
			{9'd50, 8'd77}: color_data = 12'h023;
			{9'd50, 8'd170}: color_data = 12'h000;
			{9'd50, 8'd171}: color_data = 12'h057;
			{9'd50, 8'd172}: color_data = 12'h0ae;
			{9'd50, 8'd173}: color_data = 12'h09e;
			{9'd50, 8'd174}: color_data = 12'h09e;
			{9'd50, 8'd175}: color_data = 12'h09e;
			{9'd50, 8'd176}: color_data = 12'h09e;
			{9'd50, 8'd177}: color_data = 12'h09e;
			{9'd50, 8'd178}: color_data = 12'h09e;
			{9'd50, 8'd179}: color_data = 12'h07b;
			{9'd50, 8'd180}: color_data = 12'h012;
			{9'd50, 8'd222}: color_data = 12'h310;
			{9'd50, 8'd223}: color_data = 12'he40;
			{9'd50, 8'd224}: color_data = 12'hc10;
			{9'd50, 8'd225}: color_data = 12'h900;
			{9'd50, 8'd226}: color_data = 12'h100;
			{9'd50, 8'd227}: color_data = 12'h600;
			{9'd50, 8'd228}: color_data = 12'ha00;
			{9'd50, 8'd229}: color_data = 12'ha00;
			{9'd50, 8'd230}: color_data = 12'h300;
			{9'd50, 8'd231}: color_data = 12'h720;
			{9'd50, 8'd232}: color_data = 12'hf30;
			{9'd50, 8'd233}: color_data = 12'hc10;
			{9'd50, 8'd234}: color_data = 12'h700;
			{9'd50, 8'd235}: color_data = 12'h100;
			{9'd50, 8'd236}: color_data = 12'h800;
			{9'd50, 8'd237}: color_data = 12'ha00;
			{9'd50, 8'd238}: color_data = 12'h800;
			{9'd50, 8'd239}: color_data = 12'h100;
			{9'd51, 8'd68}: color_data = 12'h057;
			{9'd51, 8'd69}: color_data = 12'h4ef;
			{9'd51, 8'd70}: color_data = 12'h7ef;
			{9'd51, 8'd71}: color_data = 12'h0cf;
			{9'd51, 8'd72}: color_data = 12'h0cf;
			{9'd51, 8'd73}: color_data = 12'h0df;
			{9'd51, 8'd74}: color_data = 12'h0bd;
			{9'd51, 8'd75}: color_data = 12'h068;
			{9'd51, 8'd76}: color_data = 12'h09c;
			{9'd51, 8'd77}: color_data = 12'h034;
			{9'd51, 8'd170}: color_data = 12'h000;
			{9'd51, 8'd171}: color_data = 12'h069;
			{9'd51, 8'd172}: color_data = 12'h6ef;
			{9'd51, 8'd173}: color_data = 12'h6ef;
			{9'd51, 8'd174}: color_data = 12'h0cf;
			{9'd51, 8'd175}: color_data = 12'h0cf;
			{9'd51, 8'd176}: color_data = 12'h0df;
			{9'd51, 8'd177}: color_data = 12'h0ac;
			{9'd51, 8'd178}: color_data = 12'h079;
			{9'd51, 8'd179}: color_data = 12'h09c;
			{9'd51, 8'd180}: color_data = 12'h023;
			{9'd51, 8'd222}: color_data = 12'h300;
			{9'd51, 8'd223}: color_data = 12'hc30;
			{9'd51, 8'd224}: color_data = 12'hd30;
			{9'd51, 8'd225}: color_data = 12'h800;
			{9'd51, 8'd226}: color_data = 12'h100;
			{9'd51, 8'd227}: color_data = 12'h600;
			{9'd51, 8'd228}: color_data = 12'ha00;
			{9'd51, 8'd229}: color_data = 12'h900;
			{9'd51, 8'd230}: color_data = 12'h300;
			{9'd51, 8'd231}: color_data = 12'h510;
			{9'd51, 8'd232}: color_data = 12'he40;
			{9'd51, 8'd233}: color_data = 12'hc20;
			{9'd51, 8'd234}: color_data = 12'h500;
			{9'd51, 8'd235}: color_data = 12'h100;
			{9'd51, 8'd236}: color_data = 12'h800;
			{9'd51, 8'd237}: color_data = 12'h900;
			{9'd51, 8'd238}: color_data = 12'h900;
			{9'd51, 8'd239}: color_data = 12'h600;
			{9'd52, 8'd68}: color_data = 12'h047;
			{9'd52, 8'd69}: color_data = 12'h6df;
			{9'd52, 8'd70}: color_data = 12'heff;
			{9'd52, 8'd71}: color_data = 12'h6df;
			{9'd52, 8'd72}: color_data = 12'h0bf;
			{9'd52, 8'd73}: color_data = 12'h0bf;
			{9'd52, 8'd74}: color_data = 12'h056;
			{9'd52, 8'd75}: color_data = 12'h012;
			{9'd52, 8'd76}: color_data = 12'h08b;
			{9'd52, 8'd77}: color_data = 12'h034;
			{9'd52, 8'd170}: color_data = 12'h000;
			{9'd52, 8'd171}: color_data = 12'h068;
			{9'd52, 8'd172}: color_data = 12'h8ef;
			{9'd52, 8'd173}: color_data = 12'hdff;
			{9'd52, 8'd174}: color_data = 12'h4cf;
			{9'd52, 8'd175}: color_data = 12'h0bf;
			{9'd52, 8'd176}: color_data = 12'h0ae;
			{9'd52, 8'd177}: color_data = 12'h035;
			{9'd52, 8'd178}: color_data = 12'h023;
			{9'd52, 8'd179}: color_data = 12'h08c;
			{9'd52, 8'd180}: color_data = 12'h023;
			{9'd52, 8'd222}: color_data = 12'h000;
			{9'd52, 8'd223}: color_data = 12'h200;
			{9'd52, 8'd224}: color_data = 12'h200;
			{9'd52, 8'd225}: color_data = 12'h100;
			{9'd52, 8'd226}: color_data = 12'h000;
			{9'd52, 8'd227}: color_data = 12'h700;
			{9'd52, 8'd228}: color_data = 12'ha00;
			{9'd52, 8'd229}: color_data = 12'h900;
			{9'd52, 8'd230}: color_data = 12'h400;
			{9'd52, 8'd231}: color_data = 12'h000;
			{9'd52, 8'd232}: color_data = 12'h200;
			{9'd52, 8'd233}: color_data = 12'h200;
			{9'd52, 8'd234}: color_data = 12'h000;
			{9'd52, 8'd235}: color_data = 12'h100;
			{9'd52, 8'd236}: color_data = 12'h800;
			{9'd52, 8'd237}: color_data = 12'ha00;
			{9'd52, 8'd238}: color_data = 12'h900;
			{9'd52, 8'd239}: color_data = 12'h500;
			{9'd53, 8'd68}: color_data = 12'h047;
			{9'd53, 8'd69}: color_data = 12'h6df;
			{9'd53, 8'd70}: color_data = 12'hfff;
			{9'd53, 8'd71}: color_data = 12'hdff;
			{9'd53, 8'd72}: color_data = 12'h5df;
			{9'd53, 8'd73}: color_data = 12'h068;
			{9'd53, 8'd74}: color_data = 12'h000;
			{9'd53, 8'd75}: color_data = 12'h012;
			{9'd53, 8'd76}: color_data = 12'h08c;
			{9'd53, 8'd77}: color_data = 12'h034;
			{9'd53, 8'd170}: color_data = 12'h000;
			{9'd53, 8'd171}: color_data = 12'h068;
			{9'd53, 8'd172}: color_data = 12'h8ef;
			{9'd53, 8'd173}: color_data = 12'hfff;
			{9'd53, 8'd174}: color_data = 12'hcff;
			{9'd53, 8'd175}: color_data = 12'h4ce;
			{9'd53, 8'd176}: color_data = 12'h057;
			{9'd53, 8'd177}: color_data = 12'h000;
			{9'd53, 8'd178}: color_data = 12'h023;
			{9'd53, 8'd179}: color_data = 12'h08c;
			{9'd53, 8'd180}: color_data = 12'h023;
			{9'd53, 8'd222}: color_data = 12'h100;
			{9'd53, 8'd223}: color_data = 12'h500;
			{9'd53, 8'd224}: color_data = 12'h600;
			{9'd53, 8'd225}: color_data = 12'h500;
			{9'd53, 8'd226}: color_data = 12'h100;
			{9'd53, 8'd227}: color_data = 12'ha20;
			{9'd53, 8'd228}: color_data = 12'hb10;
			{9'd53, 8'd229}: color_data = 12'h900;
			{9'd53, 8'd230}: color_data = 12'h400;
			{9'd53, 8'd231}: color_data = 12'h200;
			{9'd53, 8'd232}: color_data = 12'h600;
			{9'd53, 8'd233}: color_data = 12'h600;
			{9'd53, 8'd234}: color_data = 12'h400;
			{9'd53, 8'd235}: color_data = 12'h200;
			{9'd53, 8'd236}: color_data = 12'hc20;
			{9'd53, 8'd237}: color_data = 12'ha00;
			{9'd53, 8'd238}: color_data = 12'h800;
			{9'd53, 8'd239}: color_data = 12'h000;
			{9'd54, 8'd68}: color_data = 12'h047;
			{9'd54, 8'd69}: color_data = 12'h6df;
			{9'd54, 8'd70}: color_data = 12'hfff;
			{9'd54, 8'd71}: color_data = 12'hfff;
			{9'd54, 8'd72}: color_data = 12'h9aa;
			{9'd54, 8'd73}: color_data = 12'h011;
			{9'd54, 8'd75}: color_data = 12'h012;
			{9'd54, 8'd76}: color_data = 12'h08c;
			{9'd54, 8'd77}: color_data = 12'h034;
			{9'd54, 8'd170}: color_data = 12'h000;
			{9'd54, 8'd171}: color_data = 12'h068;
			{9'd54, 8'd172}: color_data = 12'h7ef;
			{9'd54, 8'd173}: color_data = 12'hfff;
			{9'd54, 8'd174}: color_data = 12'hfff;
			{9'd54, 8'd175}: color_data = 12'h899;
			{9'd54, 8'd176}: color_data = 12'h001;
			{9'd54, 8'd178}: color_data = 12'h024;
			{9'd54, 8'd179}: color_data = 12'h08c;
			{9'd54, 8'd180}: color_data = 12'h023;
			{9'd54, 8'd222}: color_data = 12'h200;
			{9'd54, 8'd223}: color_data = 12'h900;
			{9'd54, 8'd224}: color_data = 12'ha00;
			{9'd54, 8'd225}: color_data = 12'h900;
			{9'd54, 8'd226}: color_data = 12'h200;
			{9'd54, 8'd227}: color_data = 12'hb30;
			{9'd54, 8'd228}: color_data = 12'hc10;
			{9'd54, 8'd229}: color_data = 12'h900;
			{9'd54, 8'd230}: color_data = 12'h300;
			{9'd54, 8'd231}: color_data = 12'h300;
			{9'd54, 8'd232}: color_data = 12'ha00;
			{9'd54, 8'd233}: color_data = 12'ha00;
			{9'd54, 8'd234}: color_data = 12'h600;
			{9'd54, 8'd235}: color_data = 12'h310;
			{9'd54, 8'd236}: color_data = 12'he30;
			{9'd54, 8'd237}: color_data = 12'ha00;
			{9'd54, 8'd238}: color_data = 12'h700;
			{9'd54, 8'd239}: color_data = 12'h000;
			{9'd55, 8'd68}: color_data = 12'h047;
			{9'd55, 8'd69}: color_data = 12'h6df;
			{9'd55, 8'd70}: color_data = 12'hfff;
			{9'd55, 8'd71}: color_data = 12'hcbb;
			{9'd55, 8'd72}: color_data = 12'h323;
			{9'd55, 8'd73}: color_data = 12'h002;
			{9'd55, 8'd74}: color_data = 12'h000;
			{9'd55, 8'd75}: color_data = 12'h012;
			{9'd55, 8'd76}: color_data = 12'h08c;
			{9'd55, 8'd77}: color_data = 12'h034;
			{9'd55, 8'd170}: color_data = 12'h000;
			{9'd55, 8'd171}: color_data = 12'h068;
			{9'd55, 8'd172}: color_data = 12'h8ef;
			{9'd55, 8'd173}: color_data = 12'hfff;
			{9'd55, 8'd174}: color_data = 12'haaa;
			{9'd55, 8'd175}: color_data = 12'h213;
			{9'd55, 8'd176}: color_data = 12'h002;
			{9'd55, 8'd178}: color_data = 12'h023;
			{9'd55, 8'd179}: color_data = 12'h08c;
			{9'd55, 8'd180}: color_data = 12'h023;
			{9'd55, 8'd222}: color_data = 12'h200;
			{9'd55, 8'd223}: color_data = 12'h900;
			{9'd55, 8'd224}: color_data = 12'ha00;
			{9'd55, 8'd225}: color_data = 12'h800;
			{9'd55, 8'd226}: color_data = 12'h100;
			{9'd55, 8'd227}: color_data = 12'hb30;
			{9'd55, 8'd228}: color_data = 12'he30;
			{9'd55, 8'd229}: color_data = 12'hb00;
			{9'd55, 8'd230}: color_data = 12'h400;
			{9'd55, 8'd231}: color_data = 12'h300;
			{9'd55, 8'd232}: color_data = 12'h900;
			{9'd55, 8'd233}: color_data = 12'ha00;
			{9'd55, 8'd234}: color_data = 12'h600;
			{9'd55, 8'd235}: color_data = 12'h310;
			{9'd55, 8'd236}: color_data = 12'he40;
			{9'd55, 8'd237}: color_data = 12'hd20;
			{9'd55, 8'd238}: color_data = 12'h800;
			{9'd55, 8'd239}: color_data = 12'h000;
			{9'd56, 8'd68}: color_data = 12'h047;
			{9'd56, 8'd69}: color_data = 12'h6ef;
			{9'd56, 8'd70}: color_data = 12'hddc;
			{9'd56, 8'd71}: color_data = 12'h434;
			{9'd56, 8'd72}: color_data = 12'h003;
			{9'd56, 8'd73}: color_data = 12'h005;
			{9'd56, 8'd74}: color_data = 12'h002;
			{9'd56, 8'd75}: color_data = 12'h012;
			{9'd56, 8'd76}: color_data = 12'h08c;
			{9'd56, 8'd77}: color_data = 12'h034;
			{9'd56, 8'd170}: color_data = 12'h000;
			{9'd56, 8'd171}: color_data = 12'h068;
			{9'd56, 8'd172}: color_data = 12'h8ff;
			{9'd56, 8'd173}: color_data = 12'hcbb;
			{9'd56, 8'd174}: color_data = 12'h223;
			{9'd56, 8'd175}: color_data = 12'h003;
			{9'd56, 8'd176}: color_data = 12'h005;
			{9'd56, 8'd177}: color_data = 12'h002;
			{9'd56, 8'd178}: color_data = 12'h023;
			{9'd56, 8'd179}: color_data = 12'h09c;
			{9'd56, 8'd180}: color_data = 12'h023;
			{9'd56, 8'd222}: color_data = 12'h100;
			{9'd56, 8'd223}: color_data = 12'h800;
			{9'd56, 8'd224}: color_data = 12'ha00;
			{9'd56, 8'd225}: color_data = 12'h800;
			{9'd56, 8'd226}: color_data = 12'h100;
			{9'd56, 8'd227}: color_data = 12'h920;
			{9'd56, 8'd228}: color_data = 12'hd40;
			{9'd56, 8'd229}: color_data = 12'ha10;
			{9'd56, 8'd230}: color_data = 12'h200;
			{9'd56, 8'd231}: color_data = 12'h300;
			{9'd56, 8'd232}: color_data = 12'h900;
			{9'd56, 8'd233}: color_data = 12'ha00;
			{9'd56, 8'd234}: color_data = 12'h600;
			{9'd56, 8'd235}: color_data = 12'h200;
			{9'd56, 8'd236}: color_data = 12'hb30;
			{9'd56, 8'd237}: color_data = 12'hd30;
			{9'd56, 8'd238}: color_data = 12'h700;
			{9'd56, 8'd239}: color_data = 12'h000;
			{9'd57, 8'd68}: color_data = 12'h057;
			{9'd57, 8'd69}: color_data = 12'h3bd;
			{9'd57, 8'd70}: color_data = 12'h555;
			{9'd57, 8'd71}: color_data = 12'h002;
			{9'd57, 8'd72}: color_data = 12'h005;
			{9'd57, 8'd73}: color_data = 12'h005;
			{9'd57, 8'd74}: color_data = 12'h004;
			{9'd57, 8'd75}: color_data = 12'h025;
			{9'd57, 8'd76}: color_data = 12'h09c;
			{9'd57, 8'd77}: color_data = 12'h034;
			{9'd57, 8'd170}: color_data = 12'h000;
			{9'd57, 8'd171}: color_data = 12'h079;
			{9'd57, 8'd172}: color_data = 12'h4bd;
			{9'd57, 8'd173}: color_data = 12'h444;
			{9'd57, 8'd174}: color_data = 12'h002;
			{9'd57, 8'd175}: color_data = 12'h005;
			{9'd57, 8'd176}: color_data = 12'h005;
			{9'd57, 8'd177}: color_data = 12'h004;
			{9'd57, 8'd178}: color_data = 12'h036;
			{9'd57, 8'd179}: color_data = 12'h09c;
			{9'd57, 8'd180}: color_data = 12'h023;
			{9'd57, 8'd222}: color_data = 12'h200;
			{9'd57, 8'd223}: color_data = 12'h900;
			{9'd57, 8'd224}: color_data = 12'ha00;
			{9'd57, 8'd225}: color_data = 12'h900;
			{9'd57, 8'd226}: color_data = 12'h100;
			{9'd57, 8'd227}: color_data = 12'h100;
			{9'd57, 8'd228}: color_data = 12'h200;
			{9'd57, 8'd229}: color_data = 12'h100;
			{9'd57, 8'd230}: color_data = 12'h000;
			{9'd57, 8'd231}: color_data = 12'h400;
			{9'd57, 8'd232}: color_data = 12'ha00;
			{9'd57, 8'd233}: color_data = 12'ha00;
			{9'd57, 8'd234}: color_data = 12'h700;
			{9'd57, 8'd235}: color_data = 12'h000;
			{9'd57, 8'd236}: color_data = 12'h100;
			{9'd57, 8'd237}: color_data = 12'h200;
			{9'd57, 8'd238}: color_data = 12'h100;
			{9'd58, 8'd68}: color_data = 12'h035;
			{9'd58, 8'd69}: color_data = 12'h047;
			{9'd58, 8'd70}: color_data = 12'h001;
			{9'd58, 8'd71}: color_data = 12'h004;
			{9'd58, 8'd72}: color_data = 12'h004;
			{9'd58, 8'd73}: color_data = 12'h004;
			{9'd58, 8'd74}: color_data = 12'h004;
			{9'd58, 8'd75}: color_data = 12'h015;
			{9'd58, 8'd76}: color_data = 12'h059;
			{9'd58, 8'd77}: color_data = 12'h023;
			{9'd58, 8'd170}: color_data = 12'h000;
			{9'd58, 8'd171}: color_data = 12'h047;
			{9'd58, 8'd172}: color_data = 12'h036;
			{9'd58, 8'd173}: color_data = 12'h001;
			{9'd58, 8'd174}: color_data = 12'h004;
			{9'd58, 8'd175}: color_data = 12'h004;
			{9'd58, 8'd176}: color_data = 12'h004;
			{9'd58, 8'd177}: color_data = 12'h004;
			{9'd58, 8'd178}: color_data = 12'h016;
			{9'd58, 8'd179}: color_data = 12'h059;
			{9'd58, 8'd180}: color_data = 12'h012;
			{9'd58, 8'd222}: color_data = 12'h300;
			{9'd58, 8'd223}: color_data = 12'hd20;
			{9'd58, 8'd224}: color_data = 12'ha00;
			{9'd58, 8'd225}: color_data = 12'h800;
			{9'd58, 8'd226}: color_data = 12'h100;
			{9'd58, 8'd227}: color_data = 12'h400;
			{9'd58, 8'd228}: color_data = 12'h600;
			{9'd58, 8'd229}: color_data = 12'h600;
			{9'd58, 8'd230}: color_data = 12'h200;
			{9'd58, 8'd231}: color_data = 12'h610;
			{9'd58, 8'd232}: color_data = 12'hd20;
			{9'd58, 8'd233}: color_data = 12'h900;
			{9'd58, 8'd234}: color_data = 12'h600;
			{9'd58, 8'd235}: color_data = 12'h100;
			{9'd58, 8'd236}: color_data = 12'h500;
			{9'd58, 8'd237}: color_data = 12'h600;
			{9'd58, 8'd238}: color_data = 12'h500;
			{9'd58, 8'd239}: color_data = 12'h000;
			{9'd59, 8'd68}: color_data = 12'h013;
			{9'd59, 8'd69}: color_data = 12'h027;
			{9'd59, 8'd70}: color_data = 12'h016;
			{9'd59, 8'd71}: color_data = 12'h027;
			{9'd59, 8'd72}: color_data = 12'h027;
			{9'd59, 8'd73}: color_data = 12'h017;
			{9'd59, 8'd74}: color_data = 12'h027;
			{9'd59, 8'd75}: color_data = 12'h028;
			{9'd59, 8'd76}: color_data = 12'h027;
			{9'd59, 8'd77}: color_data = 12'h001;
			{9'd59, 8'd170}: color_data = 12'h000;
			{9'd59, 8'd171}: color_data = 12'h014;
			{9'd59, 8'd172}: color_data = 12'h027;
			{9'd59, 8'd173}: color_data = 12'h016;
			{9'd59, 8'd174}: color_data = 12'h027;
			{9'd59, 8'd175}: color_data = 12'h027;
			{9'd59, 8'd176}: color_data = 12'h017;
			{9'd59, 8'd177}: color_data = 12'h027;
			{9'd59, 8'd178}: color_data = 12'h028;
			{9'd59, 8'd179}: color_data = 12'h026;
			{9'd59, 8'd180}: color_data = 12'h001;
			{9'd59, 8'd222}: color_data = 12'h310;
			{9'd59, 8'd223}: color_data = 12'he30;
			{9'd59, 8'd224}: color_data = 12'ha00;
			{9'd59, 8'd225}: color_data = 12'h800;
			{9'd59, 8'd226}: color_data = 12'h100;
			{9'd59, 8'd227}: color_data = 12'h700;
			{9'd59, 8'd228}: color_data = 12'ha00;
			{9'd59, 8'd229}: color_data = 12'ha00;
			{9'd59, 8'd230}: color_data = 12'h300;
			{9'd59, 8'd231}: color_data = 12'h720;
			{9'd59, 8'd232}: color_data = 12'he30;
			{9'd59, 8'd233}: color_data = 12'h900;
			{9'd59, 8'd234}: color_data = 12'h600;
			{9'd59, 8'd235}: color_data = 12'h100;
			{9'd59, 8'd236}: color_data = 12'h900;
			{9'd59, 8'd237}: color_data = 12'ha00;
			{9'd59, 8'd238}: color_data = 12'h800;
			{9'd59, 8'd239}: color_data = 12'h000;
			{9'd60, 8'd68}: color_data = 12'h035;
			{9'd60, 8'd69}: color_data = 12'h09e;
			{9'd60, 8'd70}: color_data = 12'h09e;
			{9'd60, 8'd71}: color_data = 12'h09e;
			{9'd60, 8'd72}: color_data = 12'h09e;
			{9'd60, 8'd73}: color_data = 12'h09e;
			{9'd60, 8'd74}: color_data = 12'h09e;
			{9'd60, 8'd75}: color_data = 12'h09e;
			{9'd60, 8'd76}: color_data = 12'h08c;
			{9'd60, 8'd77}: color_data = 12'h023;
			{9'd60, 8'd170}: color_data = 12'h000;
			{9'd60, 8'd171}: color_data = 12'h057;
			{9'd60, 8'd172}: color_data = 12'h0ae;
			{9'd60, 8'd173}: color_data = 12'h09e;
			{9'd60, 8'd174}: color_data = 12'h09e;
			{9'd60, 8'd175}: color_data = 12'h09e;
			{9'd60, 8'd176}: color_data = 12'h09e;
			{9'd60, 8'd177}: color_data = 12'h09e;
			{9'd60, 8'd178}: color_data = 12'h09e;
			{9'd60, 8'd179}: color_data = 12'h07b;
			{9'd60, 8'd180}: color_data = 12'h012;
			{9'd60, 8'd222}: color_data = 12'h310;
			{9'd60, 8'd223}: color_data = 12'hf40;
			{9'd60, 8'd224}: color_data = 12'hd20;
			{9'd60, 8'd225}: color_data = 12'h900;
			{9'd60, 8'd226}: color_data = 12'h100;
			{9'd60, 8'd227}: color_data = 12'h600;
			{9'd60, 8'd228}: color_data = 12'ha00;
			{9'd60, 8'd229}: color_data = 12'h900;
			{9'd60, 8'd230}: color_data = 12'h300;
			{9'd60, 8'd231}: color_data = 12'h720;
			{9'd60, 8'd232}: color_data = 12'hf40;
			{9'd60, 8'd233}: color_data = 12'hc10;
			{9'd60, 8'd234}: color_data = 12'h700;
			{9'd60, 8'd235}: color_data = 12'h100;
			{9'd60, 8'd236}: color_data = 12'h800;
			{9'd60, 8'd237}: color_data = 12'ha00;
			{9'd60, 8'd238}: color_data = 12'h800;
			{9'd60, 8'd239}: color_data = 12'h100;
			{9'd61, 8'd68}: color_data = 12'h057;
			{9'd61, 8'd69}: color_data = 12'h4ef;
			{9'd61, 8'd70}: color_data = 12'h7ef;
			{9'd61, 8'd71}: color_data = 12'h0cf;
			{9'd61, 8'd72}: color_data = 12'h0cf;
			{9'd61, 8'd73}: color_data = 12'h0df;
			{9'd61, 8'd74}: color_data = 12'h0bd;
			{9'd61, 8'd75}: color_data = 12'h068;
			{9'd61, 8'd76}: color_data = 12'h09c;
			{9'd61, 8'd77}: color_data = 12'h034;
			{9'd61, 8'd170}: color_data = 12'h000;
			{9'd61, 8'd171}: color_data = 12'h069;
			{9'd61, 8'd172}: color_data = 12'h6ef;
			{9'd61, 8'd173}: color_data = 12'h6ef;
			{9'd61, 8'd174}: color_data = 12'h0cf;
			{9'd61, 8'd175}: color_data = 12'h0cf;
			{9'd61, 8'd176}: color_data = 12'h0df;
			{9'd61, 8'd177}: color_data = 12'h0ac;
			{9'd61, 8'd178}: color_data = 12'h079;
			{9'd61, 8'd179}: color_data = 12'h09c;
			{9'd61, 8'd180}: color_data = 12'h023;
			{9'd61, 8'd222}: color_data = 12'h200;
			{9'd61, 8'd223}: color_data = 12'hb30;
			{9'd61, 8'd224}: color_data = 12'hc30;
			{9'd61, 8'd225}: color_data = 12'h700;
			{9'd61, 8'd226}: color_data = 12'h100;
			{9'd61, 8'd227}: color_data = 12'h600;
			{9'd61, 8'd228}: color_data = 12'ha00;
			{9'd61, 8'd229}: color_data = 12'h900;
			{9'd61, 8'd230}: color_data = 12'h300;
			{9'd61, 8'd231}: color_data = 12'h410;
			{9'd61, 8'd232}: color_data = 12'hc40;
			{9'd61, 8'd233}: color_data = 12'hb20;
			{9'd61, 8'd234}: color_data = 12'h500;
			{9'd61, 8'd235}: color_data = 12'h100;
			{9'd61, 8'd236}: color_data = 12'h800;
			{9'd61, 8'd237}: color_data = 12'ha00;
			{9'd61, 8'd238}: color_data = 12'h800;
			{9'd61, 8'd239}: color_data = 12'h100;
			{9'd62, 8'd68}: color_data = 12'h047;
			{9'd62, 8'd69}: color_data = 12'h6df;
			{9'd62, 8'd70}: color_data = 12'heff;
			{9'd62, 8'd71}: color_data = 12'h6df;
			{9'd62, 8'd72}: color_data = 12'h0bf;
			{9'd62, 8'd73}: color_data = 12'h0bf;
			{9'd62, 8'd74}: color_data = 12'h056;
			{9'd62, 8'd75}: color_data = 12'h012;
			{9'd62, 8'd76}: color_data = 12'h08b;
			{9'd62, 8'd77}: color_data = 12'h034;
			{9'd62, 8'd170}: color_data = 12'h000;
			{9'd62, 8'd171}: color_data = 12'h068;
			{9'd62, 8'd172}: color_data = 12'h8ef;
			{9'd62, 8'd173}: color_data = 12'hdff;
			{9'd62, 8'd174}: color_data = 12'h4cf;
			{9'd62, 8'd175}: color_data = 12'h0bf;
			{9'd62, 8'd176}: color_data = 12'h0ae;
			{9'd62, 8'd177}: color_data = 12'h045;
			{9'd62, 8'd178}: color_data = 12'h023;
			{9'd62, 8'd179}: color_data = 12'h08c;
			{9'd62, 8'd180}: color_data = 12'h023;
			{9'd62, 8'd222}: color_data = 12'h000;
			{9'd62, 8'd223}: color_data = 12'h100;
			{9'd62, 8'd224}: color_data = 12'h100;
			{9'd62, 8'd225}: color_data = 12'h100;
			{9'd62, 8'd226}: color_data = 12'h000;
			{9'd62, 8'd227}: color_data = 12'h700;
			{9'd62, 8'd228}: color_data = 12'ha00;
			{9'd62, 8'd229}: color_data = 12'h900;
			{9'd62, 8'd230}: color_data = 12'h400;
			{9'd62, 8'd231}: color_data = 12'h000;
			{9'd62, 8'd232}: color_data = 12'h100;
			{9'd62, 8'd233}: color_data = 12'h100;
			{9'd62, 8'd234}: color_data = 12'h000;
			{9'd62, 8'd235}: color_data = 12'h100;
			{9'd62, 8'd236}: color_data = 12'h900;
			{9'd62, 8'd237}: color_data = 12'ha00;
			{9'd62, 8'd238}: color_data = 12'h800;
			{9'd62, 8'd239}: color_data = 12'h100;
			{9'd63, 8'd68}: color_data = 12'h047;
			{9'd63, 8'd69}: color_data = 12'h6df;
			{9'd63, 8'd70}: color_data = 12'hfff;
			{9'd63, 8'd71}: color_data = 12'hdff;
			{9'd63, 8'd72}: color_data = 12'h5df;
			{9'd63, 8'd73}: color_data = 12'h068;
			{9'd63, 8'd74}: color_data = 12'h000;
			{9'd63, 8'd75}: color_data = 12'h012;
			{9'd63, 8'd76}: color_data = 12'h08c;
			{9'd63, 8'd77}: color_data = 12'h034;
			{9'd63, 8'd170}: color_data = 12'h000;
			{9'd63, 8'd171}: color_data = 12'h068;
			{9'd63, 8'd172}: color_data = 12'h8ef;
			{9'd63, 8'd173}: color_data = 12'hfff;
			{9'd63, 8'd174}: color_data = 12'hcff;
			{9'd63, 8'd175}: color_data = 12'h4ce;
			{9'd63, 8'd176}: color_data = 12'h057;
			{9'd63, 8'd177}: color_data = 12'h000;
			{9'd63, 8'd178}: color_data = 12'h023;
			{9'd63, 8'd179}: color_data = 12'h08c;
			{9'd63, 8'd180}: color_data = 12'h023;
			{9'd63, 8'd222}: color_data = 12'h100;
			{9'd63, 8'd223}: color_data = 12'h600;
			{9'd63, 8'd224}: color_data = 12'h700;
			{9'd63, 8'd225}: color_data = 12'h600;
			{9'd63, 8'd226}: color_data = 12'h100;
			{9'd63, 8'd227}: color_data = 12'ha20;
			{9'd63, 8'd228}: color_data = 12'hc10;
			{9'd63, 8'd229}: color_data = 12'h900;
			{9'd63, 8'd230}: color_data = 12'h400;
			{9'd63, 8'd231}: color_data = 12'h200;
			{9'd63, 8'd232}: color_data = 12'h700;
			{9'd63, 8'd233}: color_data = 12'h700;
			{9'd63, 8'd234}: color_data = 12'h400;
			{9'd63, 8'd235}: color_data = 12'h200;
			{9'd63, 8'd236}: color_data = 12'hd20;
			{9'd63, 8'd237}: color_data = 12'ha00;
			{9'd63, 8'd238}: color_data = 12'h800;
			{9'd63, 8'd239}: color_data = 12'h100;
			{9'd64, 8'd68}: color_data = 12'h047;
			{9'd64, 8'd69}: color_data = 12'h6df;
			{9'd64, 8'd70}: color_data = 12'hfff;
			{9'd64, 8'd71}: color_data = 12'hfff;
			{9'd64, 8'd72}: color_data = 12'h9aa;
			{9'd64, 8'd73}: color_data = 12'h011;
			{9'd64, 8'd75}: color_data = 12'h012;
			{9'd64, 8'd76}: color_data = 12'h08c;
			{9'd64, 8'd77}: color_data = 12'h034;
			{9'd64, 8'd170}: color_data = 12'h000;
			{9'd64, 8'd171}: color_data = 12'h068;
			{9'd64, 8'd172}: color_data = 12'h7ef;
			{9'd64, 8'd173}: color_data = 12'hfff;
			{9'd64, 8'd174}: color_data = 12'hfff;
			{9'd64, 8'd175}: color_data = 12'h899;
			{9'd64, 8'd176}: color_data = 12'h001;
			{9'd64, 8'd178}: color_data = 12'h024;
			{9'd64, 8'd179}: color_data = 12'h08c;
			{9'd64, 8'd180}: color_data = 12'h023;
			{9'd64, 8'd222}: color_data = 12'h200;
			{9'd64, 8'd223}: color_data = 12'h900;
			{9'd64, 8'd224}: color_data = 12'ha00;
			{9'd64, 8'd225}: color_data = 12'h900;
			{9'd64, 8'd226}: color_data = 12'h200;
			{9'd64, 8'd227}: color_data = 12'hb30;
			{9'd64, 8'd228}: color_data = 12'hc10;
			{9'd64, 8'd229}: color_data = 12'h900;
			{9'd64, 8'd230}: color_data = 12'h300;
			{9'd64, 8'd231}: color_data = 12'h300;
			{9'd64, 8'd232}: color_data = 12'ha00;
			{9'd64, 8'd233}: color_data = 12'ha00;
			{9'd64, 8'd234}: color_data = 12'h600;
			{9'd64, 8'd235}: color_data = 12'h310;
			{9'd64, 8'd236}: color_data = 12'he30;
			{9'd64, 8'd237}: color_data = 12'ha00;
			{9'd64, 8'd238}: color_data = 12'h800;
			{9'd64, 8'd239}: color_data = 12'h000;
			{9'd65, 8'd68}: color_data = 12'h047;
			{9'd65, 8'd69}: color_data = 12'h6df;
			{9'd65, 8'd70}: color_data = 12'hfff;
			{9'd65, 8'd71}: color_data = 12'hcbb;
			{9'd65, 8'd72}: color_data = 12'h323;
			{9'd65, 8'd73}: color_data = 12'h002;
			{9'd65, 8'd74}: color_data = 12'h000;
			{9'd65, 8'd75}: color_data = 12'h012;
			{9'd65, 8'd76}: color_data = 12'h08c;
			{9'd65, 8'd77}: color_data = 12'h034;
			{9'd65, 8'd170}: color_data = 12'h000;
			{9'd65, 8'd171}: color_data = 12'h068;
			{9'd65, 8'd172}: color_data = 12'h8ef;
			{9'd65, 8'd173}: color_data = 12'hfff;
			{9'd65, 8'd174}: color_data = 12'haaa;
			{9'd65, 8'd175}: color_data = 12'h213;
			{9'd65, 8'd176}: color_data = 12'h002;
			{9'd65, 8'd178}: color_data = 12'h023;
			{9'd65, 8'd179}: color_data = 12'h08c;
			{9'd65, 8'd180}: color_data = 12'h023;
			{9'd65, 8'd222}: color_data = 12'h200;
			{9'd65, 8'd223}: color_data = 12'h900;
			{9'd65, 8'd224}: color_data = 12'ha00;
			{9'd65, 8'd225}: color_data = 12'h800;
			{9'd65, 8'd226}: color_data = 12'h100;
			{9'd65, 8'd227}: color_data = 12'hb30;
			{9'd65, 8'd228}: color_data = 12'hf30;
			{9'd65, 8'd229}: color_data = 12'hb00;
			{9'd65, 8'd230}: color_data = 12'h400;
			{9'd65, 8'd231}: color_data = 12'h300;
			{9'd65, 8'd232}: color_data = 12'h900;
			{9'd65, 8'd233}: color_data = 12'ha00;
			{9'd65, 8'd234}: color_data = 12'h600;
			{9'd65, 8'd235}: color_data = 12'h310;
			{9'd65, 8'd236}: color_data = 12'he40;
			{9'd65, 8'd237}: color_data = 12'he20;
			{9'd65, 8'd238}: color_data = 12'h900;
			{9'd65, 8'd239}: color_data = 12'h000;
			{9'd66, 8'd68}: color_data = 12'h047;
			{9'd66, 8'd69}: color_data = 12'h6ef;
			{9'd66, 8'd70}: color_data = 12'hdcc;
			{9'd66, 8'd71}: color_data = 12'h434;
			{9'd66, 8'd72}: color_data = 12'h003;
			{9'd66, 8'd73}: color_data = 12'h005;
			{9'd66, 8'd74}: color_data = 12'h002;
			{9'd66, 8'd75}: color_data = 12'h012;
			{9'd66, 8'd76}: color_data = 12'h08c;
			{9'd66, 8'd77}: color_data = 12'h034;
			{9'd66, 8'd170}: color_data = 12'h000;
			{9'd66, 8'd171}: color_data = 12'h068;
			{9'd66, 8'd172}: color_data = 12'h8ff;
			{9'd66, 8'd173}: color_data = 12'hcbb;
			{9'd66, 8'd174}: color_data = 12'h323;
			{9'd66, 8'd175}: color_data = 12'h003;
			{9'd66, 8'd176}: color_data = 12'h005;
			{9'd66, 8'd177}: color_data = 12'h002;
			{9'd66, 8'd178}: color_data = 12'h023;
			{9'd66, 8'd179}: color_data = 12'h09c;
			{9'd66, 8'd180}: color_data = 12'h023;
			{9'd66, 8'd222}: color_data = 12'h100;
			{9'd66, 8'd223}: color_data = 12'h800;
			{9'd66, 8'd224}: color_data = 12'ha00;
			{9'd66, 8'd225}: color_data = 12'h800;
			{9'd66, 8'd226}: color_data = 12'h100;
			{9'd66, 8'd227}: color_data = 12'h820;
			{9'd66, 8'd228}: color_data = 12'hc30;
			{9'd66, 8'd229}: color_data = 12'h910;
			{9'd66, 8'd230}: color_data = 12'h200;
			{9'd66, 8'd231}: color_data = 12'h300;
			{9'd66, 8'd232}: color_data = 12'h900;
			{9'd66, 8'd233}: color_data = 12'ha00;
			{9'd66, 8'd234}: color_data = 12'h600;
			{9'd66, 8'd235}: color_data = 12'h200;
			{9'd66, 8'd236}: color_data = 12'ha30;
			{9'd66, 8'd237}: color_data = 12'hc30;
			{9'd66, 8'd238}: color_data = 12'h700;
			{9'd66, 8'd239}: color_data = 12'h000;
			{9'd67, 8'd68}: color_data = 12'h057;
			{9'd67, 8'd69}: color_data = 12'h3bd;
			{9'd67, 8'd70}: color_data = 12'h555;
			{9'd67, 8'd71}: color_data = 12'h002;
			{9'd67, 8'd72}: color_data = 12'h005;
			{9'd67, 8'd73}: color_data = 12'h005;
			{9'd67, 8'd74}: color_data = 12'h004;
			{9'd67, 8'd75}: color_data = 12'h025;
			{9'd67, 8'd76}: color_data = 12'h09c;
			{9'd67, 8'd77}: color_data = 12'h034;
			{9'd67, 8'd170}: color_data = 12'h000;
			{9'd67, 8'd171}: color_data = 12'h079;
			{9'd67, 8'd172}: color_data = 12'h4bd;
			{9'd67, 8'd173}: color_data = 12'h444;
			{9'd67, 8'd174}: color_data = 12'h002;
			{9'd67, 8'd175}: color_data = 12'h005;
			{9'd67, 8'd176}: color_data = 12'h005;
			{9'd67, 8'd177}: color_data = 12'h004;
			{9'd67, 8'd178}: color_data = 12'h036;
			{9'd67, 8'd179}: color_data = 12'h09c;
			{9'd67, 8'd180}: color_data = 12'h023;
			{9'd67, 8'd222}: color_data = 12'h200;
			{9'd67, 8'd223}: color_data = 12'h900;
			{9'd67, 8'd224}: color_data = 12'ha00;
			{9'd67, 8'd225}: color_data = 12'h900;
			{9'd67, 8'd226}: color_data = 12'h100;
			{9'd67, 8'd227}: color_data = 12'h000;
			{9'd67, 8'd228}: color_data = 12'h100;
			{9'd67, 8'd229}: color_data = 12'h100;
			{9'd67, 8'd230}: color_data = 12'h000;
			{9'd67, 8'd231}: color_data = 12'h400;
			{9'd67, 8'd232}: color_data = 12'ha00;
			{9'd67, 8'd233}: color_data = 12'ha00;
			{9'd67, 8'd234}: color_data = 12'h700;
			{9'd67, 8'd235}: color_data = 12'h000;
			{9'd67, 8'd236}: color_data = 12'h100;
			{9'd67, 8'd237}: color_data = 12'h100;
			{9'd67, 8'd238}: color_data = 12'h100;
			{9'd67, 8'd239}: color_data = 12'h100;
			{9'd68, 8'd68}: color_data = 12'h035;
			{9'd68, 8'd69}: color_data = 12'h047;
			{9'd68, 8'd70}: color_data = 12'h001;
			{9'd68, 8'd71}: color_data = 12'h004;
			{9'd68, 8'd72}: color_data = 12'h004;
			{9'd68, 8'd73}: color_data = 12'h004;
			{9'd68, 8'd74}: color_data = 12'h004;
			{9'd68, 8'd75}: color_data = 12'h015;
			{9'd68, 8'd76}: color_data = 12'h059;
			{9'd68, 8'd77}: color_data = 12'h023;
			{9'd68, 8'd170}: color_data = 12'h000;
			{9'd68, 8'd171}: color_data = 12'h047;
			{9'd68, 8'd172}: color_data = 12'h036;
			{9'd68, 8'd173}: color_data = 12'h001;
			{9'd68, 8'd174}: color_data = 12'h004;
			{9'd68, 8'd175}: color_data = 12'h004;
			{9'd68, 8'd176}: color_data = 12'h004;
			{9'd68, 8'd177}: color_data = 12'h004;
			{9'd68, 8'd178}: color_data = 12'h016;
			{9'd68, 8'd179}: color_data = 12'h059;
			{9'd68, 8'd180}: color_data = 12'h012;
			{9'd68, 8'd222}: color_data = 12'h310;
			{9'd68, 8'd223}: color_data = 12'hd30;
			{9'd68, 8'd224}: color_data = 12'ha00;
			{9'd68, 8'd225}: color_data = 12'h800;
			{9'd68, 8'd226}: color_data = 12'h100;
			{9'd68, 8'd227}: color_data = 12'h400;
			{9'd68, 8'd228}: color_data = 12'h700;
			{9'd68, 8'd229}: color_data = 12'h700;
			{9'd68, 8'd230}: color_data = 12'h200;
			{9'd68, 8'd231}: color_data = 12'h610;
			{9'd68, 8'd232}: color_data = 12'hd20;
			{9'd68, 8'd233}: color_data = 12'h900;
			{9'd68, 8'd234}: color_data = 12'h600;
			{9'd68, 8'd235}: color_data = 12'h100;
			{9'd68, 8'd236}: color_data = 12'h600;
			{9'd68, 8'd237}: color_data = 12'h700;
			{9'd68, 8'd238}: color_data = 12'h700;
			{9'd68, 8'd239}: color_data = 12'h100;
			{9'd69, 8'd68}: color_data = 12'h013;
			{9'd69, 8'd69}: color_data = 12'h027;
			{9'd69, 8'd70}: color_data = 12'h016;
			{9'd69, 8'd71}: color_data = 12'h027;
			{9'd69, 8'd72}: color_data = 12'h027;
			{9'd69, 8'd73}: color_data = 12'h027;
			{9'd69, 8'd74}: color_data = 12'h027;
			{9'd69, 8'd75}: color_data = 12'h028;
			{9'd69, 8'd76}: color_data = 12'h027;
			{9'd69, 8'd77}: color_data = 12'h001;
			{9'd69, 8'd119}: color_data = 12'h000;
			{9'd69, 8'd120}: color_data = 12'h012;
			{9'd69, 8'd121}: color_data = 12'h023;
			{9'd69, 8'd122}: color_data = 12'h022;
			{9'd69, 8'd123}: color_data = 12'h022;
			{9'd69, 8'd124}: color_data = 12'h022;
			{9'd69, 8'd125}: color_data = 12'h022;
			{9'd69, 8'd126}: color_data = 12'h023;
			{9'd69, 8'd127}: color_data = 12'h023;
			{9'd69, 8'd128}: color_data = 12'h011;
			{9'd69, 8'd170}: color_data = 12'h000;
			{9'd69, 8'd171}: color_data = 12'h014;
			{9'd69, 8'd172}: color_data = 12'h027;
			{9'd69, 8'd173}: color_data = 12'h016;
			{9'd69, 8'd174}: color_data = 12'h027;
			{9'd69, 8'd175}: color_data = 12'h027;
			{9'd69, 8'd176}: color_data = 12'h027;
			{9'd69, 8'd177}: color_data = 12'h027;
			{9'd69, 8'd178}: color_data = 12'h028;
			{9'd69, 8'd179}: color_data = 12'h026;
			{9'd69, 8'd180}: color_data = 12'h001;
			{9'd69, 8'd222}: color_data = 12'h310;
			{9'd69, 8'd223}: color_data = 12'he30;
			{9'd69, 8'd224}: color_data = 12'ha00;
			{9'd69, 8'd225}: color_data = 12'h800;
			{9'd69, 8'd226}: color_data = 12'h100;
			{9'd69, 8'd227}: color_data = 12'h600;
			{9'd69, 8'd228}: color_data = 12'ha00;
			{9'd69, 8'd229}: color_data = 12'ha00;
			{9'd69, 8'd230}: color_data = 12'h300;
			{9'd69, 8'd231}: color_data = 12'h720;
			{9'd69, 8'd232}: color_data = 12'he30;
			{9'd69, 8'd233}: color_data = 12'h900;
			{9'd69, 8'd234}: color_data = 12'h600;
			{9'd69, 8'd235}: color_data = 12'h100;
			{9'd69, 8'd236}: color_data = 12'h900;
			{9'd69, 8'd237}: color_data = 12'ha00;
			{9'd69, 8'd238}: color_data = 12'h900;
			{9'd69, 8'd239}: color_data = 12'h100;
			{9'd70, 8'd68}: color_data = 12'h036;
			{9'd70, 8'd69}: color_data = 12'h09e;
			{9'd70, 8'd70}: color_data = 12'h09e;
			{9'd70, 8'd71}: color_data = 12'h09e;
			{9'd70, 8'd72}: color_data = 12'h09e;
			{9'd70, 8'd73}: color_data = 12'h09e;
			{9'd70, 8'd74}: color_data = 12'h09e;
			{9'd70, 8'd75}: color_data = 12'h09e;
			{9'd70, 8'd76}: color_data = 12'h08c;
			{9'd70, 8'd77}: color_data = 12'h023;
			{9'd70, 8'd119}: color_data = 12'h012;
			{9'd70, 8'd120}: color_data = 12'h08b;
			{9'd70, 8'd121}: color_data = 12'h0ad;
			{9'd70, 8'd122}: color_data = 12'h09d;
			{9'd70, 8'd123}: color_data = 12'h09d;
			{9'd70, 8'd124}: color_data = 12'h09d;
			{9'd70, 8'd125}: color_data = 12'h09d;
			{9'd70, 8'd126}: color_data = 12'h09d;
			{9'd70, 8'd127}: color_data = 12'h09d;
			{9'd70, 8'd128}: color_data = 12'h057;
			{9'd70, 8'd129}: color_data = 12'h000;
			{9'd70, 8'd170}: color_data = 12'h000;
			{9'd70, 8'd171}: color_data = 12'h057;
			{9'd70, 8'd172}: color_data = 12'h0ae;
			{9'd70, 8'd173}: color_data = 12'h09e;
			{9'd70, 8'd174}: color_data = 12'h09e;
			{9'd70, 8'd175}: color_data = 12'h09e;
			{9'd70, 8'd176}: color_data = 12'h09e;
			{9'd70, 8'd177}: color_data = 12'h09e;
			{9'd70, 8'd178}: color_data = 12'h09e;
			{9'd70, 8'd179}: color_data = 12'h07b;
			{9'd70, 8'd180}: color_data = 12'h012;
			{9'd70, 8'd222}: color_data = 12'h310;
			{9'd70, 8'd223}: color_data = 12'hf40;
			{9'd70, 8'd224}: color_data = 12'he20;
			{9'd70, 8'd225}: color_data = 12'h900;
			{9'd70, 8'd226}: color_data = 12'h100;
			{9'd70, 8'd227}: color_data = 12'h600;
			{9'd70, 8'd228}: color_data = 12'ha00;
			{9'd70, 8'd229}: color_data = 12'h900;
			{9'd70, 8'd230}: color_data = 12'h300;
			{9'd70, 8'd231}: color_data = 12'h720;
			{9'd70, 8'd232}: color_data = 12'hf40;
			{9'd70, 8'd233}: color_data = 12'hd10;
			{9'd70, 8'd234}: color_data = 12'h700;
			{9'd70, 8'd235}: color_data = 12'h100;
			{9'd70, 8'd236}: color_data = 12'h800;
			{9'd70, 8'd237}: color_data = 12'ha00;
			{9'd70, 8'd238}: color_data = 12'h800;
			{9'd70, 8'd239}: color_data = 12'h100;
			{9'd71, 8'd68}: color_data = 12'h057;
			{9'd71, 8'd69}: color_data = 12'h4ef;
			{9'd71, 8'd70}: color_data = 12'h7ef;
			{9'd71, 8'd71}: color_data = 12'h0cf;
			{9'd71, 8'd72}: color_data = 12'h0cf;
			{9'd71, 8'd73}: color_data = 12'h0df;
			{9'd71, 8'd74}: color_data = 12'h0bd;
			{9'd71, 8'd75}: color_data = 12'h068;
			{9'd71, 8'd76}: color_data = 12'h09c;
			{9'd71, 8'd77}: color_data = 12'h034;
			{9'd71, 8'd119}: color_data = 12'h012;
			{9'd71, 8'd120}: color_data = 12'h1bd;
			{9'd71, 8'd121}: color_data = 12'h8ff;
			{9'd71, 8'd122}: color_data = 12'h3df;
			{9'd71, 8'd123}: color_data = 12'h0cf;
			{9'd71, 8'd124}: color_data = 12'h0cf;
			{9'd71, 8'd125}: color_data = 12'h0cf;
			{9'd71, 8'd126}: color_data = 12'h07a;
			{9'd71, 8'd127}: color_data = 12'h08b;
			{9'd71, 8'd128}: color_data = 12'h079;
			{9'd71, 8'd129}: color_data = 12'h000;
			{9'd71, 8'd170}: color_data = 12'h000;
			{9'd71, 8'd171}: color_data = 12'h069;
			{9'd71, 8'd172}: color_data = 12'h6ef;
			{9'd71, 8'd173}: color_data = 12'h6ef;
			{9'd71, 8'd174}: color_data = 12'h0cf;
			{9'd71, 8'd175}: color_data = 12'h0cf;
			{9'd71, 8'd176}: color_data = 12'h0df;
			{9'd71, 8'd177}: color_data = 12'h0ac;
			{9'd71, 8'd178}: color_data = 12'h079;
			{9'd71, 8'd179}: color_data = 12'h09c;
			{9'd71, 8'd180}: color_data = 12'h023;
			{9'd71, 8'd222}: color_data = 12'h200;
			{9'd71, 8'd223}: color_data = 12'ha30;
			{9'd71, 8'd224}: color_data = 12'hb30;
			{9'd71, 8'd225}: color_data = 12'h600;
			{9'd71, 8'd226}: color_data = 12'h100;
			{9'd71, 8'd227}: color_data = 12'h600;
			{9'd71, 8'd228}: color_data = 12'h900;
			{9'd71, 8'd229}: color_data = 12'h900;
			{9'd71, 8'd230}: color_data = 12'h300;
			{9'd71, 8'd231}: color_data = 12'h410;
			{9'd71, 8'd232}: color_data = 12'hb30;
			{9'd71, 8'd233}: color_data = 12'ha20;
			{9'd71, 8'd234}: color_data = 12'h400;
			{9'd71, 8'd235}: color_data = 12'h100;
			{9'd71, 8'd236}: color_data = 12'h800;
			{9'd71, 8'd237}: color_data = 12'ha00;
			{9'd71, 8'd238}: color_data = 12'h800;
			{9'd71, 8'd239}: color_data = 12'h100;
			{9'd72, 8'd68}: color_data = 12'h047;
			{9'd72, 8'd69}: color_data = 12'h6df;
			{9'd72, 8'd70}: color_data = 12'heff;
			{9'd72, 8'd71}: color_data = 12'h6df;
			{9'd72, 8'd72}: color_data = 12'h0bf;
			{9'd72, 8'd73}: color_data = 12'h0bf;
			{9'd72, 8'd74}: color_data = 12'h056;
			{9'd72, 8'd75}: color_data = 12'h012;
			{9'd72, 8'd76}: color_data = 12'h08b;
			{9'd72, 8'd77}: color_data = 12'h034;
			{9'd72, 8'd119}: color_data = 12'h012;
			{9'd72, 8'd120}: color_data = 12'h2ad;
			{9'd72, 8'd121}: color_data = 12'hdff;
			{9'd72, 8'd122}: color_data = 12'haef;
			{9'd72, 8'd123}: color_data = 12'h1bf;
			{9'd72, 8'd124}: color_data = 12'h0cf;
			{9'd72, 8'd125}: color_data = 12'h08b;
			{9'd72, 8'd126}: color_data = 12'h012;
			{9'd72, 8'd127}: color_data = 12'h068;
			{9'd72, 8'd128}: color_data = 12'h079;
			{9'd72, 8'd129}: color_data = 12'h000;
			{9'd72, 8'd170}: color_data = 12'h000;
			{9'd72, 8'd171}: color_data = 12'h068;
			{9'd72, 8'd172}: color_data = 12'h8ef;
			{9'd72, 8'd173}: color_data = 12'hdff;
			{9'd72, 8'd174}: color_data = 12'h4cf;
			{9'd72, 8'd175}: color_data = 12'h0bf;
			{9'd72, 8'd176}: color_data = 12'h0ae;
			{9'd72, 8'd177}: color_data = 12'h035;
			{9'd72, 8'd178}: color_data = 12'h023;
			{9'd72, 8'd179}: color_data = 12'h08c;
			{9'd72, 8'd180}: color_data = 12'h023;
			{9'd72, 8'd222}: color_data = 12'h000;
			{9'd72, 8'd223}: color_data = 12'h100;
			{9'd72, 8'd224}: color_data = 12'h100;
			{9'd72, 8'd225}: color_data = 12'h100;
			{9'd72, 8'd226}: color_data = 12'h000;
			{9'd72, 8'd227}: color_data = 12'h700;
			{9'd72, 8'd228}: color_data = 12'ha00;
			{9'd72, 8'd229}: color_data = 12'h900;
			{9'd72, 8'd230}: color_data = 12'h400;
			{9'd72, 8'd231}: color_data = 12'h000;
			{9'd72, 8'd232}: color_data = 12'h100;
			{9'd72, 8'd233}: color_data = 12'h100;
			{9'd72, 8'd234}: color_data = 12'h000;
			{9'd72, 8'd235}: color_data = 12'h100;
			{9'd72, 8'd236}: color_data = 12'h900;
			{9'd72, 8'd237}: color_data = 12'ha00;
			{9'd72, 8'd238}: color_data = 12'h800;
			{9'd72, 8'd239}: color_data = 12'h100;
			{9'd73, 8'd68}: color_data = 12'h047;
			{9'd73, 8'd69}: color_data = 12'h6df;
			{9'd73, 8'd70}: color_data = 12'hfff;
			{9'd73, 8'd71}: color_data = 12'hdff;
			{9'd73, 8'd72}: color_data = 12'h5df;
			{9'd73, 8'd73}: color_data = 12'h068;
			{9'd73, 8'd74}: color_data = 12'h000;
			{9'd73, 8'd75}: color_data = 12'h012;
			{9'd73, 8'd76}: color_data = 12'h08c;
			{9'd73, 8'd77}: color_data = 12'h034;
			{9'd73, 8'd119}: color_data = 12'h012;
			{9'd73, 8'd120}: color_data = 12'h1ad;
			{9'd73, 8'd121}: color_data = 12'hdff;
			{9'd73, 8'd122}: color_data = 12'hfff;
			{9'd73, 8'd123}: color_data = 12'h8ef;
			{9'd73, 8'd124}: color_data = 12'h19c;
			{9'd73, 8'd125}: color_data = 12'h023;
			{9'd73, 8'd127}: color_data = 12'h068;
			{9'd73, 8'd128}: color_data = 12'h079;
			{9'd73, 8'd129}: color_data = 12'h000;
			{9'd73, 8'd170}: color_data = 12'h000;
			{9'd73, 8'd171}: color_data = 12'h068;
			{9'd73, 8'd172}: color_data = 12'h8ef;
			{9'd73, 8'd173}: color_data = 12'hfff;
			{9'd73, 8'd174}: color_data = 12'hcff;
			{9'd73, 8'd175}: color_data = 12'h4ce;
			{9'd73, 8'd176}: color_data = 12'h057;
			{9'd73, 8'd177}: color_data = 12'h000;
			{9'd73, 8'd178}: color_data = 12'h023;
			{9'd73, 8'd179}: color_data = 12'h08c;
			{9'd73, 8'd180}: color_data = 12'h023;
			{9'd73, 8'd222}: color_data = 12'h100;
			{9'd73, 8'd223}: color_data = 12'h700;
			{9'd73, 8'd224}: color_data = 12'h800;
			{9'd73, 8'd225}: color_data = 12'h700;
			{9'd73, 8'd226}: color_data = 12'h100;
			{9'd73, 8'd227}: color_data = 12'ha20;
			{9'd73, 8'd228}: color_data = 12'hc10;
			{9'd73, 8'd229}: color_data = 12'h900;
			{9'd73, 8'd230}: color_data = 12'h400;
			{9'd73, 8'd231}: color_data = 12'h200;
			{9'd73, 8'd232}: color_data = 12'h800;
			{9'd73, 8'd233}: color_data = 12'h800;
			{9'd73, 8'd234}: color_data = 12'h500;
			{9'd73, 8'd235}: color_data = 12'h200;
			{9'd73, 8'd236}: color_data = 12'hd30;
			{9'd73, 8'd237}: color_data = 12'ha00;
			{9'd73, 8'd238}: color_data = 12'h800;
			{9'd73, 8'd239}: color_data = 12'h100;
			{9'd74, 8'd68}: color_data = 12'h047;
			{9'd74, 8'd69}: color_data = 12'h6df;
			{9'd74, 8'd70}: color_data = 12'hfff;
			{9'd74, 8'd71}: color_data = 12'hfff;
			{9'd74, 8'd72}: color_data = 12'h9aa;
			{9'd74, 8'd73}: color_data = 12'h011;
			{9'd74, 8'd75}: color_data = 12'h012;
			{9'd74, 8'd76}: color_data = 12'h08c;
			{9'd74, 8'd77}: color_data = 12'h034;
			{9'd74, 8'd119}: color_data = 12'h012;
			{9'd74, 8'd120}: color_data = 12'h1ad;
			{9'd74, 8'd121}: color_data = 12'hcff;
			{9'd74, 8'd122}: color_data = 12'hfff;
			{9'd74, 8'd123}: color_data = 12'hddd;
			{9'd74, 8'd124}: color_data = 12'h345;
			{9'd74, 8'd126}: color_data = 12'h000;
			{9'd74, 8'd127}: color_data = 12'h068;
			{9'd74, 8'd128}: color_data = 12'h079;
			{9'd74, 8'd129}: color_data = 12'h000;
			{9'd74, 8'd170}: color_data = 12'h000;
			{9'd74, 8'd171}: color_data = 12'h068;
			{9'd74, 8'd172}: color_data = 12'h7ef;
			{9'd74, 8'd173}: color_data = 12'hfff;
			{9'd74, 8'd174}: color_data = 12'hfff;
			{9'd74, 8'd175}: color_data = 12'h899;
			{9'd74, 8'd176}: color_data = 12'h001;
			{9'd74, 8'd178}: color_data = 12'h024;
			{9'd74, 8'd179}: color_data = 12'h08c;
			{9'd74, 8'd180}: color_data = 12'h023;
			{9'd74, 8'd222}: color_data = 12'h200;
			{9'd74, 8'd223}: color_data = 12'h900;
			{9'd74, 8'd224}: color_data = 12'ha00;
			{9'd74, 8'd225}: color_data = 12'h900;
			{9'd74, 8'd226}: color_data = 12'h200;
			{9'd74, 8'd227}: color_data = 12'hb30;
			{9'd74, 8'd228}: color_data = 12'hc10;
			{9'd74, 8'd229}: color_data = 12'h900;
			{9'd74, 8'd230}: color_data = 12'h300;
			{9'd74, 8'd231}: color_data = 12'h300;
			{9'd74, 8'd232}: color_data = 12'ha00;
			{9'd74, 8'd233}: color_data = 12'ha00;
			{9'd74, 8'd234}: color_data = 12'h600;
			{9'd74, 8'd235}: color_data = 12'h310;
			{9'd74, 8'd236}: color_data = 12'he30;
			{9'd74, 8'd237}: color_data = 12'ha00;
			{9'd74, 8'd238}: color_data = 12'h800;
			{9'd74, 8'd239}: color_data = 12'h000;
			{9'd75, 8'd68}: color_data = 12'h047;
			{9'd75, 8'd69}: color_data = 12'h6df;
			{9'd75, 8'd70}: color_data = 12'hfff;
			{9'd75, 8'd71}: color_data = 12'hcbb;
			{9'd75, 8'd72}: color_data = 12'h323;
			{9'd75, 8'd73}: color_data = 12'h002;
			{9'd75, 8'd74}: color_data = 12'h000;
			{9'd75, 8'd75}: color_data = 12'h012;
			{9'd75, 8'd76}: color_data = 12'h08c;
			{9'd75, 8'd77}: color_data = 12'h034;
			{9'd75, 8'd119}: color_data = 12'h012;
			{9'd75, 8'd120}: color_data = 12'h1ad;
			{9'd75, 8'd121}: color_data = 12'hdff;
			{9'd75, 8'd122}: color_data = 12'hfee;
			{9'd75, 8'd123}: color_data = 12'h666;
			{9'd75, 8'd124}: color_data = 12'h002;
			{9'd75, 8'd125}: color_data = 12'h001;
			{9'd75, 8'd126}: color_data = 12'h000;
			{9'd75, 8'd127}: color_data = 12'h068;
			{9'd75, 8'd128}: color_data = 12'h079;
			{9'd75, 8'd129}: color_data = 12'h000;
			{9'd75, 8'd170}: color_data = 12'h000;
			{9'd75, 8'd171}: color_data = 12'h068;
			{9'd75, 8'd172}: color_data = 12'h8ef;
			{9'd75, 8'd173}: color_data = 12'hfff;
			{9'd75, 8'd174}: color_data = 12'haaa;
			{9'd75, 8'd175}: color_data = 12'h213;
			{9'd75, 8'd176}: color_data = 12'h002;
			{9'd75, 8'd178}: color_data = 12'h023;
			{9'd75, 8'd179}: color_data = 12'h08c;
			{9'd75, 8'd180}: color_data = 12'h023;
			{9'd75, 8'd222}: color_data = 12'h200;
			{9'd75, 8'd223}: color_data = 12'h900;
			{9'd75, 8'd224}: color_data = 12'ha00;
			{9'd75, 8'd225}: color_data = 12'h800;
			{9'd75, 8'd226}: color_data = 12'h100;
			{9'd75, 8'd227}: color_data = 12'hb30;
			{9'd75, 8'd228}: color_data = 12'hf30;
			{9'd75, 8'd229}: color_data = 12'hc00;
			{9'd75, 8'd230}: color_data = 12'h300;
			{9'd75, 8'd231}: color_data = 12'h300;
			{9'd75, 8'd232}: color_data = 12'h900;
			{9'd75, 8'd233}: color_data = 12'ha00;
			{9'd75, 8'd234}: color_data = 12'h600;
			{9'd75, 8'd235}: color_data = 12'h310;
			{9'd75, 8'd236}: color_data = 12'he40;
			{9'd75, 8'd237}: color_data = 12'he20;
			{9'd75, 8'd238}: color_data = 12'h900;
			{9'd75, 8'd239}: color_data = 12'h000;
			{9'd76, 8'd68}: color_data = 12'h047;
			{9'd76, 8'd69}: color_data = 12'h6ef;
			{9'd76, 8'd70}: color_data = 12'hddc;
			{9'd76, 8'd71}: color_data = 12'h434;
			{9'd76, 8'd72}: color_data = 12'h003;
			{9'd76, 8'd73}: color_data = 12'h005;
			{9'd76, 8'd74}: color_data = 12'h002;
			{9'd76, 8'd75}: color_data = 12'h012;
			{9'd76, 8'd76}: color_data = 12'h08c;
			{9'd76, 8'd77}: color_data = 12'h034;
			{9'd76, 8'd119}: color_data = 12'h012;
			{9'd76, 8'd120}: color_data = 12'h2ad;
			{9'd76, 8'd121}: color_data = 12'hcff;
			{9'd76, 8'd122}: color_data = 12'h877;
			{9'd76, 8'd123}: color_data = 12'h002;
			{9'd76, 8'd124}: color_data = 12'h004;
			{9'd76, 8'd125}: color_data = 12'h004;
			{9'd76, 8'd126}: color_data = 12'h000;
			{9'd76, 8'd127}: color_data = 12'h068;
			{9'd76, 8'd128}: color_data = 12'h079;
			{9'd76, 8'd129}: color_data = 12'h000;
			{9'd76, 8'd170}: color_data = 12'h000;
			{9'd76, 8'd171}: color_data = 12'h068;
			{9'd76, 8'd172}: color_data = 12'h8ff;
			{9'd76, 8'd173}: color_data = 12'hcbb;
			{9'd76, 8'd174}: color_data = 12'h323;
			{9'd76, 8'd175}: color_data = 12'h003;
			{9'd76, 8'd176}: color_data = 12'h005;
			{9'd76, 8'd177}: color_data = 12'h002;
			{9'd76, 8'd178}: color_data = 12'h023;
			{9'd76, 8'd179}: color_data = 12'h09c;
			{9'd76, 8'd180}: color_data = 12'h023;
			{9'd76, 8'd222}: color_data = 12'h100;
			{9'd76, 8'd223}: color_data = 12'h800;
			{9'd76, 8'd224}: color_data = 12'ha00;
			{9'd76, 8'd225}: color_data = 12'h800;
			{9'd76, 8'd226}: color_data = 12'h100;
			{9'd76, 8'd227}: color_data = 12'h720;
			{9'd76, 8'd228}: color_data = 12'hb30;
			{9'd76, 8'd229}: color_data = 12'h810;
			{9'd76, 8'd230}: color_data = 12'h100;
			{9'd76, 8'd231}: color_data = 12'h300;
			{9'd76, 8'd232}: color_data = 12'h900;
			{9'd76, 8'd233}: color_data = 12'ha00;
			{9'd76, 8'd234}: color_data = 12'h600;
			{9'd76, 8'd235}: color_data = 12'h100;
			{9'd76, 8'd236}: color_data = 12'h930;
			{9'd76, 8'd237}: color_data = 12'ha30;
			{9'd76, 8'd238}: color_data = 12'h600;
			{9'd76, 8'd239}: color_data = 12'h000;
			{9'd77, 8'd68}: color_data = 12'h057;
			{9'd77, 8'd69}: color_data = 12'h3bd;
			{9'd77, 8'd70}: color_data = 12'h555;
			{9'd77, 8'd71}: color_data = 12'h002;
			{9'd77, 8'd72}: color_data = 12'h005;
			{9'd77, 8'd73}: color_data = 12'h005;
			{9'd77, 8'd74}: color_data = 12'h004;
			{9'd77, 8'd75}: color_data = 12'h025;
			{9'd77, 8'd76}: color_data = 12'h09c;
			{9'd77, 8'd77}: color_data = 12'h034;
			{9'd77, 8'd119}: color_data = 12'h022;
			{9'd77, 8'd120}: color_data = 12'h1ad;
			{9'd77, 8'd121}: color_data = 12'h689;
			{9'd77, 8'd122}: color_data = 12'h212;
			{9'd77, 8'd123}: color_data = 12'h004;
			{9'd77, 8'd124}: color_data = 12'h005;
			{9'd77, 8'd125}: color_data = 12'h005;
			{9'd77, 8'd126}: color_data = 12'h003;
			{9'd77, 8'd127}: color_data = 12'h06a;
			{9'd77, 8'd128}: color_data = 12'h079;
			{9'd77, 8'd129}: color_data = 12'h000;
			{9'd77, 8'd170}: color_data = 12'h000;
			{9'd77, 8'd171}: color_data = 12'h079;
			{9'd77, 8'd172}: color_data = 12'h4bd;
			{9'd77, 8'd173}: color_data = 12'h444;
			{9'd77, 8'd174}: color_data = 12'h002;
			{9'd77, 8'd175}: color_data = 12'h005;
			{9'd77, 8'd176}: color_data = 12'h005;
			{9'd77, 8'd177}: color_data = 12'h004;
			{9'd77, 8'd178}: color_data = 12'h036;
			{9'd77, 8'd179}: color_data = 12'h09c;
			{9'd77, 8'd180}: color_data = 12'h023;
			{9'd77, 8'd222}: color_data = 12'h200;
			{9'd77, 8'd223}: color_data = 12'h900;
			{9'd77, 8'd224}: color_data = 12'ha00;
			{9'd77, 8'd225}: color_data = 12'h900;
			{9'd77, 8'd226}: color_data = 12'h100;
			{9'd77, 8'd227}: color_data = 12'h000;
			{9'd77, 8'd228}: color_data = 12'h100;
			{9'd77, 8'd229}: color_data = 12'h100;
			{9'd77, 8'd230}: color_data = 12'h000;
			{9'd77, 8'd231}: color_data = 12'h400;
			{9'd77, 8'd232}: color_data = 12'ha00;
			{9'd77, 8'd233}: color_data = 12'ha00;
			{9'd77, 8'd234}: color_data = 12'h700;
			{9'd77, 8'd235}: color_data = 12'h000;
			{9'd77, 8'd236}: color_data = 12'h100;
			{9'd77, 8'd237}: color_data = 12'h100;
			{9'd77, 8'd238}: color_data = 12'h100;
			{9'd77, 8'd239}: color_data = 12'h100;
			{9'd78, 8'd68}: color_data = 12'h035;
			{9'd78, 8'd69}: color_data = 12'h047;
			{9'd78, 8'd70}: color_data = 12'h001;
			{9'd78, 8'd71}: color_data = 12'h004;
			{9'd78, 8'd72}: color_data = 12'h004;
			{9'd78, 8'd73}: color_data = 12'h004;
			{9'd78, 8'd74}: color_data = 12'h004;
			{9'd78, 8'd75}: color_data = 12'h015;
			{9'd78, 8'd76}: color_data = 12'h059;
			{9'd78, 8'd77}: color_data = 12'h023;
			{9'd78, 8'd119}: color_data = 12'h012;
			{9'd78, 8'd120}: color_data = 12'h059;
			{9'd78, 8'd121}: color_data = 12'h013;
			{9'd78, 8'd122}: color_data = 12'h002;
			{9'd78, 8'd123}: color_data = 12'h004;
			{9'd78, 8'd124}: color_data = 12'h004;
			{9'd78, 8'd125}: color_data = 12'h004;
			{9'd78, 8'd126}: color_data = 12'h004;
			{9'd78, 8'd127}: color_data = 12'h039;
			{9'd78, 8'd128}: color_data = 12'h047;
			{9'd78, 8'd129}: color_data = 12'h000;
			{9'd78, 8'd170}: color_data = 12'h000;
			{9'd78, 8'd171}: color_data = 12'h047;
			{9'd78, 8'd172}: color_data = 12'h036;
			{9'd78, 8'd173}: color_data = 12'h001;
			{9'd78, 8'd174}: color_data = 12'h004;
			{9'd78, 8'd175}: color_data = 12'h004;
			{9'd78, 8'd176}: color_data = 12'h004;
			{9'd78, 8'd177}: color_data = 12'h004;
			{9'd78, 8'd178}: color_data = 12'h016;
			{9'd78, 8'd179}: color_data = 12'h059;
			{9'd78, 8'd180}: color_data = 12'h012;
			{9'd78, 8'd222}: color_data = 12'h310;
			{9'd78, 8'd223}: color_data = 12'hd30;
			{9'd78, 8'd224}: color_data = 12'ha00;
			{9'd78, 8'd225}: color_data = 12'h800;
			{9'd78, 8'd226}: color_data = 12'h100;
			{9'd78, 8'd227}: color_data = 12'h500;
			{9'd78, 8'd228}: color_data = 12'h800;
			{9'd78, 8'd229}: color_data = 12'h800;
			{9'd78, 8'd230}: color_data = 12'h300;
			{9'd78, 8'd231}: color_data = 12'h620;
			{9'd78, 8'd232}: color_data = 12'hd20;
			{9'd78, 8'd233}: color_data = 12'h900;
			{9'd78, 8'd234}: color_data = 12'h600;
			{9'd78, 8'd235}: color_data = 12'h100;
			{9'd78, 8'd236}: color_data = 12'h700;
			{9'd78, 8'd237}: color_data = 12'h800;
			{9'd78, 8'd238}: color_data = 12'h700;
			{9'd78, 8'd239}: color_data = 12'h100;
			{9'd79, 8'd68}: color_data = 12'h013;
			{9'd79, 8'd69}: color_data = 12'h027;
			{9'd79, 8'd70}: color_data = 12'h016;
			{9'd79, 8'd71}: color_data = 12'h027;
			{9'd79, 8'd72}: color_data = 12'h027;
			{9'd79, 8'd73}: color_data = 12'h017;
			{9'd79, 8'd74}: color_data = 12'h027;
			{9'd79, 8'd75}: color_data = 12'h028;
			{9'd79, 8'd76}: color_data = 12'h027;
			{9'd79, 8'd77}: color_data = 12'h001;
			{9'd79, 8'd119}: color_data = 12'h001;
			{9'd79, 8'd120}: color_data = 12'h016;
			{9'd79, 8'd121}: color_data = 12'h017;
			{9'd79, 8'd122}: color_data = 12'h016;
			{9'd79, 8'd123}: color_data = 12'h027;
			{9'd79, 8'd124}: color_data = 12'h027;
			{9'd79, 8'd125}: color_data = 12'h027;
			{9'd79, 8'd126}: color_data = 12'h027;
			{9'd79, 8'd127}: color_data = 12'h028;
			{9'd79, 8'd128}: color_data = 12'h014;
			{9'd79, 8'd129}: color_data = 12'h000;
			{9'd79, 8'd170}: color_data = 12'h000;
			{9'd79, 8'd171}: color_data = 12'h014;
			{9'd79, 8'd172}: color_data = 12'h027;
			{9'd79, 8'd173}: color_data = 12'h016;
			{9'd79, 8'd174}: color_data = 12'h027;
			{9'd79, 8'd175}: color_data = 12'h027;
			{9'd79, 8'd176}: color_data = 12'h017;
			{9'd79, 8'd177}: color_data = 12'h027;
			{9'd79, 8'd178}: color_data = 12'h028;
			{9'd79, 8'd179}: color_data = 12'h026;
			{9'd79, 8'd180}: color_data = 12'h001;
			{9'd79, 8'd222}: color_data = 12'h310;
			{9'd79, 8'd223}: color_data = 12'he30;
			{9'd79, 8'd224}: color_data = 12'ha00;
			{9'd79, 8'd225}: color_data = 12'h800;
			{9'd79, 8'd226}: color_data = 12'h100;
			{9'd79, 8'd227}: color_data = 12'h600;
			{9'd79, 8'd228}: color_data = 12'ha00;
			{9'd79, 8'd229}: color_data = 12'ha00;
			{9'd79, 8'd230}: color_data = 12'h300;
			{9'd79, 8'd231}: color_data = 12'h720;
			{9'd79, 8'd232}: color_data = 12'he30;
			{9'd79, 8'd233}: color_data = 12'h900;
			{9'd79, 8'd234}: color_data = 12'h600;
			{9'd79, 8'd235}: color_data = 12'h100;
			{9'd79, 8'd236}: color_data = 12'h900;
			{9'd79, 8'd237}: color_data = 12'ha00;
			{9'd79, 8'd238}: color_data = 12'h900;
			{9'd79, 8'd239}: color_data = 12'h100;
			{9'd80, 8'd68}: color_data = 12'h035;
			{9'd80, 8'd69}: color_data = 12'h09e;
			{9'd80, 8'd70}: color_data = 12'h09e;
			{9'd80, 8'd71}: color_data = 12'h09e;
			{9'd80, 8'd72}: color_data = 12'h09e;
			{9'd80, 8'd73}: color_data = 12'h09e;
			{9'd80, 8'd74}: color_data = 12'h09e;
			{9'd80, 8'd75}: color_data = 12'h09e;
			{9'd80, 8'd76}: color_data = 12'h08c;
			{9'd80, 8'd77}: color_data = 12'h023;
			{9'd80, 8'd119}: color_data = 12'h012;
			{9'd80, 8'd120}: color_data = 12'h07b;
			{9'd80, 8'd121}: color_data = 12'h0ae;
			{9'd80, 8'd122}: color_data = 12'h09e;
			{9'd80, 8'd123}: color_data = 12'h09e;
			{9'd80, 8'd124}: color_data = 12'h09e;
			{9'd80, 8'd125}: color_data = 12'h09e;
			{9'd80, 8'd126}: color_data = 12'h09e;
			{9'd80, 8'd127}: color_data = 12'h09e;
			{9'd80, 8'd128}: color_data = 12'h057;
			{9'd80, 8'd129}: color_data = 12'h000;
			{9'd80, 8'd170}: color_data = 12'h000;
			{9'd80, 8'd171}: color_data = 12'h057;
			{9'd80, 8'd172}: color_data = 12'h0ae;
			{9'd80, 8'd173}: color_data = 12'h09e;
			{9'd80, 8'd174}: color_data = 12'h09e;
			{9'd80, 8'd175}: color_data = 12'h09e;
			{9'd80, 8'd176}: color_data = 12'h09e;
			{9'd80, 8'd177}: color_data = 12'h09e;
			{9'd80, 8'd178}: color_data = 12'h09e;
			{9'd80, 8'd179}: color_data = 12'h07b;
			{9'd80, 8'd180}: color_data = 12'h012;
			{9'd80, 8'd222}: color_data = 12'h310;
			{9'd80, 8'd223}: color_data = 12'hf40;
			{9'd80, 8'd224}: color_data = 12'he20;
			{9'd80, 8'd225}: color_data = 12'ha00;
			{9'd80, 8'd226}: color_data = 12'h100;
			{9'd80, 8'd227}: color_data = 12'h600;
			{9'd80, 8'd228}: color_data = 12'ha00;
			{9'd80, 8'd229}: color_data = 12'h900;
			{9'd80, 8'd230}: color_data = 12'h300;
			{9'd80, 8'd231}: color_data = 12'h720;
			{9'd80, 8'd232}: color_data = 12'hf40;
			{9'd80, 8'd233}: color_data = 12'hd10;
			{9'd80, 8'd234}: color_data = 12'h700;
			{9'd80, 8'd235}: color_data = 12'h100;
			{9'd80, 8'd236}: color_data = 12'h800;
			{9'd80, 8'd237}: color_data = 12'ha00;
			{9'd80, 8'd238}: color_data = 12'h800;
			{9'd80, 8'd239}: color_data = 12'h100;
			{9'd81, 8'd68}: color_data = 12'h057;
			{9'd81, 8'd69}: color_data = 12'h4ef;
			{9'd81, 8'd70}: color_data = 12'h7ef;
			{9'd81, 8'd71}: color_data = 12'h0cf;
			{9'd81, 8'd72}: color_data = 12'h0cf;
			{9'd81, 8'd73}: color_data = 12'h0df;
			{9'd81, 8'd74}: color_data = 12'h0bd;
			{9'd81, 8'd75}: color_data = 12'h068;
			{9'd81, 8'd76}: color_data = 12'h09c;
			{9'd81, 8'd77}: color_data = 12'h034;
			{9'd81, 8'd119}: color_data = 12'h001;
			{9'd81, 8'd120}: color_data = 12'h1ad;
			{9'd81, 8'd121}: color_data = 12'h8ff;
			{9'd81, 8'd122}: color_data = 12'h3df;
			{9'd81, 8'd123}: color_data = 12'h0cf;
			{9'd81, 8'd124}: color_data = 12'h0cf;
			{9'd81, 8'd125}: color_data = 12'h0cf;
			{9'd81, 8'd126}: color_data = 12'h07a;
			{9'd81, 8'd127}: color_data = 12'h08b;
			{9'd81, 8'd128}: color_data = 12'h079;
			{9'd81, 8'd129}: color_data = 12'h000;
			{9'd81, 8'd170}: color_data = 12'h000;
			{9'd81, 8'd171}: color_data = 12'h069;
			{9'd81, 8'd172}: color_data = 12'h6ef;
			{9'd81, 8'd173}: color_data = 12'h6ef;
			{9'd81, 8'd174}: color_data = 12'h0cf;
			{9'd81, 8'd175}: color_data = 12'h0cf;
			{9'd81, 8'd176}: color_data = 12'h0df;
			{9'd81, 8'd177}: color_data = 12'h0ad;
			{9'd81, 8'd178}: color_data = 12'h079;
			{9'd81, 8'd179}: color_data = 12'h09c;
			{9'd81, 8'd180}: color_data = 12'h023;
			{9'd81, 8'd222}: color_data = 12'h200;
			{9'd81, 8'd223}: color_data = 12'h920;
			{9'd81, 8'd224}: color_data = 12'h920;
			{9'd81, 8'd225}: color_data = 12'h500;
			{9'd81, 8'd226}: color_data = 12'h000;
			{9'd81, 8'd227}: color_data = 12'h600;
			{9'd81, 8'd228}: color_data = 12'h900;
			{9'd81, 8'd229}: color_data = 12'h900;
			{9'd81, 8'd230}: color_data = 12'h300;
			{9'd81, 8'd231}: color_data = 12'h310;
			{9'd81, 8'd232}: color_data = 12'ha30;
			{9'd81, 8'd233}: color_data = 12'h820;
			{9'd81, 8'd234}: color_data = 12'h300;
			{9'd81, 8'd235}: color_data = 12'h100;
			{9'd81, 8'd236}: color_data = 12'h800;
			{9'd81, 8'd237}: color_data = 12'h900;
			{9'd81, 8'd238}: color_data = 12'h800;
			{9'd81, 8'd239}: color_data = 12'h100;
			{9'd82, 8'd68}: color_data = 12'h047;
			{9'd82, 8'd69}: color_data = 12'h6df;
			{9'd82, 8'd70}: color_data = 12'heff;
			{9'd82, 8'd71}: color_data = 12'h6df;
			{9'd82, 8'd72}: color_data = 12'h0bf;
			{9'd82, 8'd73}: color_data = 12'h0be;
			{9'd82, 8'd74}: color_data = 12'h056;
			{9'd82, 8'd75}: color_data = 12'h012;
			{9'd82, 8'd76}: color_data = 12'h08b;
			{9'd82, 8'd77}: color_data = 12'h034;
			{9'd82, 8'd119}: color_data = 12'h000;
			{9'd82, 8'd120}: color_data = 12'h2ac;
			{9'd82, 8'd121}: color_data = 12'hdff;
			{9'd82, 8'd122}: color_data = 12'haef;
			{9'd82, 8'd123}: color_data = 12'h1cf;
			{9'd82, 8'd124}: color_data = 12'h0cf;
			{9'd82, 8'd125}: color_data = 12'h08b;
			{9'd82, 8'd126}: color_data = 12'h012;
			{9'd82, 8'd127}: color_data = 12'h068;
			{9'd82, 8'd128}: color_data = 12'h079;
			{9'd82, 8'd129}: color_data = 12'h000;
			{9'd82, 8'd170}: color_data = 12'h000;
			{9'd82, 8'd171}: color_data = 12'h068;
			{9'd82, 8'd172}: color_data = 12'h8ef;
			{9'd82, 8'd173}: color_data = 12'hdff;
			{9'd82, 8'd174}: color_data = 12'h4cf;
			{9'd82, 8'd175}: color_data = 12'h0cf;
			{9'd82, 8'd176}: color_data = 12'h0ae;
			{9'd82, 8'd177}: color_data = 12'h035;
			{9'd82, 8'd178}: color_data = 12'h023;
			{9'd82, 8'd179}: color_data = 12'h08c;
			{9'd82, 8'd180}: color_data = 12'h023;
			{9'd82, 8'd222}: color_data = 12'h000;
			{9'd82, 8'd223}: color_data = 12'h100;
			{9'd82, 8'd224}: color_data = 12'h100;
			{9'd82, 8'd225}: color_data = 12'h100;
			{9'd82, 8'd226}: color_data = 12'h000;
			{9'd82, 8'd227}: color_data = 12'h700;
			{9'd82, 8'd228}: color_data = 12'ha00;
			{9'd82, 8'd229}: color_data = 12'h900;
			{9'd82, 8'd230}: color_data = 12'h400;
			{9'd82, 8'd231}: color_data = 12'h000;
			{9'd82, 8'd232}: color_data = 12'h100;
			{9'd82, 8'd233}: color_data = 12'h100;
			{9'd82, 8'd234}: color_data = 12'h000;
			{9'd82, 8'd235}: color_data = 12'h100;
			{9'd82, 8'd236}: color_data = 12'h900;
			{9'd82, 8'd237}: color_data = 12'ha00;
			{9'd82, 8'd238}: color_data = 12'h800;
			{9'd82, 8'd239}: color_data = 12'h100;
			{9'd83, 8'd68}: color_data = 12'h047;
			{9'd83, 8'd69}: color_data = 12'h6df;
			{9'd83, 8'd70}: color_data = 12'hfff;
			{9'd83, 8'd71}: color_data = 12'hdff;
			{9'd83, 8'd72}: color_data = 12'h5df;
			{9'd83, 8'd73}: color_data = 12'h068;
			{9'd83, 8'd74}: color_data = 12'h000;
			{9'd83, 8'd75}: color_data = 12'h012;
			{9'd83, 8'd76}: color_data = 12'h08c;
			{9'd83, 8'd77}: color_data = 12'h034;
			{9'd83, 8'd119}: color_data = 12'h000;
			{9'd83, 8'd120}: color_data = 12'h1ac;
			{9'd83, 8'd121}: color_data = 12'hdff;
			{9'd83, 8'd122}: color_data = 12'hfff;
			{9'd83, 8'd123}: color_data = 12'h8ef;
			{9'd83, 8'd124}: color_data = 12'h19c;
			{9'd83, 8'd125}: color_data = 12'h023;
			{9'd83, 8'd127}: color_data = 12'h068;
			{9'd83, 8'd128}: color_data = 12'h079;
			{9'd83, 8'd129}: color_data = 12'h000;
			{9'd83, 8'd170}: color_data = 12'h000;
			{9'd83, 8'd171}: color_data = 12'h068;
			{9'd83, 8'd172}: color_data = 12'h8ef;
			{9'd83, 8'd173}: color_data = 12'hfff;
			{9'd83, 8'd174}: color_data = 12'hcff;
			{9'd83, 8'd175}: color_data = 12'h4ce;
			{9'd83, 8'd176}: color_data = 12'h057;
			{9'd83, 8'd177}: color_data = 12'h000;
			{9'd83, 8'd178}: color_data = 12'h023;
			{9'd83, 8'd179}: color_data = 12'h08c;
			{9'd83, 8'd180}: color_data = 12'h023;
			{9'd83, 8'd222}: color_data = 12'h100;
			{9'd83, 8'd223}: color_data = 12'h800;
			{9'd83, 8'd224}: color_data = 12'h900;
			{9'd83, 8'd225}: color_data = 12'h700;
			{9'd83, 8'd226}: color_data = 12'h100;
			{9'd83, 8'd227}: color_data = 12'hb30;
			{9'd83, 8'd228}: color_data = 12'hc10;
			{9'd83, 8'd229}: color_data = 12'h900;
			{9'd83, 8'd230}: color_data = 12'h400;
			{9'd83, 8'd231}: color_data = 12'h300;
			{9'd83, 8'd232}: color_data = 12'h800;
			{9'd83, 8'd233}: color_data = 12'h900;
			{9'd83, 8'd234}: color_data = 12'h500;
			{9'd83, 8'd235}: color_data = 12'h200;
			{9'd83, 8'd236}: color_data = 12'hd30;
			{9'd83, 8'd237}: color_data = 12'ha00;
			{9'd83, 8'd238}: color_data = 12'h800;
			{9'd83, 8'd239}: color_data = 12'h100;
			{9'd84, 8'd68}: color_data = 12'h047;
			{9'd84, 8'd69}: color_data = 12'h6df;
			{9'd84, 8'd70}: color_data = 12'hfff;
			{9'd84, 8'd71}: color_data = 12'hfff;
			{9'd84, 8'd72}: color_data = 12'h9aa;
			{9'd84, 8'd73}: color_data = 12'h011;
			{9'd84, 8'd75}: color_data = 12'h012;
			{9'd84, 8'd76}: color_data = 12'h08c;
			{9'd84, 8'd77}: color_data = 12'h034;
			{9'd84, 8'd119}: color_data = 12'h000;
			{9'd84, 8'd120}: color_data = 12'h1ac;
			{9'd84, 8'd121}: color_data = 12'hcff;
			{9'd84, 8'd122}: color_data = 12'hfff;
			{9'd84, 8'd123}: color_data = 12'hddd;
			{9'd84, 8'd124}: color_data = 12'h345;
			{9'd84, 8'd126}: color_data = 12'h000;
			{9'd84, 8'd127}: color_data = 12'h068;
			{9'd84, 8'd128}: color_data = 12'h079;
			{9'd84, 8'd129}: color_data = 12'h000;
			{9'd84, 8'd170}: color_data = 12'h000;
			{9'd84, 8'd171}: color_data = 12'h068;
			{9'd84, 8'd172}: color_data = 12'h7ef;
			{9'd84, 8'd173}: color_data = 12'hfff;
			{9'd84, 8'd174}: color_data = 12'hfff;
			{9'd84, 8'd175}: color_data = 12'h899;
			{9'd84, 8'd176}: color_data = 12'h001;
			{9'd84, 8'd178}: color_data = 12'h024;
			{9'd84, 8'd179}: color_data = 12'h08c;
			{9'd84, 8'd180}: color_data = 12'h023;
			{9'd84, 8'd222}: color_data = 12'h200;
			{9'd84, 8'd223}: color_data = 12'h900;
			{9'd84, 8'd224}: color_data = 12'ha00;
			{9'd84, 8'd225}: color_data = 12'h900;
			{9'd84, 8'd226}: color_data = 12'h200;
			{9'd84, 8'd227}: color_data = 12'hb30;
			{9'd84, 8'd228}: color_data = 12'hc10;
			{9'd84, 8'd229}: color_data = 12'h900;
			{9'd84, 8'd230}: color_data = 12'h300;
			{9'd84, 8'd231}: color_data = 12'h300;
			{9'd84, 8'd232}: color_data = 12'ha00;
			{9'd84, 8'd233}: color_data = 12'ha00;
			{9'd84, 8'd234}: color_data = 12'h600;
			{9'd84, 8'd235}: color_data = 12'h310;
			{9'd84, 8'd236}: color_data = 12'he30;
			{9'd84, 8'd237}: color_data = 12'ha00;
			{9'd84, 8'd238}: color_data = 12'h800;
			{9'd84, 8'd239}: color_data = 12'h000;
			{9'd85, 8'd68}: color_data = 12'h047;
			{9'd85, 8'd69}: color_data = 12'h6df;
			{9'd85, 8'd70}: color_data = 12'hfff;
			{9'd85, 8'd71}: color_data = 12'hcbb;
			{9'd85, 8'd72}: color_data = 12'h323;
			{9'd85, 8'd73}: color_data = 12'h002;
			{9'd85, 8'd74}: color_data = 12'h000;
			{9'd85, 8'd75}: color_data = 12'h012;
			{9'd85, 8'd76}: color_data = 12'h08c;
			{9'd85, 8'd77}: color_data = 12'h034;
			{9'd85, 8'd119}: color_data = 12'h000;
			{9'd85, 8'd120}: color_data = 12'h1ac;
			{9'd85, 8'd121}: color_data = 12'hdff;
			{9'd85, 8'd122}: color_data = 12'hfee;
			{9'd85, 8'd123}: color_data = 12'h666;
			{9'd85, 8'd124}: color_data = 12'h002;
			{9'd85, 8'd125}: color_data = 12'h001;
			{9'd85, 8'd126}: color_data = 12'h000;
			{9'd85, 8'd127}: color_data = 12'h068;
			{9'd85, 8'd128}: color_data = 12'h079;
			{9'd85, 8'd129}: color_data = 12'h000;
			{9'd85, 8'd170}: color_data = 12'h000;
			{9'd85, 8'd171}: color_data = 12'h068;
			{9'd85, 8'd172}: color_data = 12'h8ef;
			{9'd85, 8'd173}: color_data = 12'hfff;
			{9'd85, 8'd174}: color_data = 12'haaa;
			{9'd85, 8'd175}: color_data = 12'h213;
			{9'd85, 8'd176}: color_data = 12'h002;
			{9'd85, 8'd178}: color_data = 12'h023;
			{9'd85, 8'd179}: color_data = 12'h08c;
			{9'd85, 8'd180}: color_data = 12'h023;
			{9'd85, 8'd222}: color_data = 12'h200;
			{9'd85, 8'd223}: color_data = 12'h900;
			{9'd85, 8'd224}: color_data = 12'ha00;
			{9'd85, 8'd225}: color_data = 12'h800;
			{9'd85, 8'd226}: color_data = 12'h100;
			{9'd85, 8'd227}: color_data = 12'hb30;
			{9'd85, 8'd228}: color_data = 12'hf40;
			{9'd85, 8'd229}: color_data = 12'hc10;
			{9'd85, 8'd230}: color_data = 12'h300;
			{9'd85, 8'd231}: color_data = 12'h300;
			{9'd85, 8'd232}: color_data = 12'h900;
			{9'd85, 8'd233}: color_data = 12'ha00;
			{9'd85, 8'd234}: color_data = 12'h600;
			{9'd85, 8'd235}: color_data = 12'h300;
			{9'd85, 8'd236}: color_data = 12'he40;
			{9'd85, 8'd237}: color_data = 12'hf30;
			{9'd85, 8'd238}: color_data = 12'h900;
			{9'd85, 8'd239}: color_data = 12'h000;
			{9'd86, 8'd68}: color_data = 12'h047;
			{9'd86, 8'd69}: color_data = 12'h6ef;
			{9'd86, 8'd70}: color_data = 12'hdcc;
			{9'd86, 8'd71}: color_data = 12'h434;
			{9'd86, 8'd72}: color_data = 12'h003;
			{9'd86, 8'd73}: color_data = 12'h005;
			{9'd86, 8'd74}: color_data = 12'h002;
			{9'd86, 8'd75}: color_data = 12'h012;
			{9'd86, 8'd76}: color_data = 12'h08c;
			{9'd86, 8'd77}: color_data = 12'h034;
			{9'd86, 8'd119}: color_data = 12'h000;
			{9'd86, 8'd120}: color_data = 12'h2ad;
			{9'd86, 8'd121}: color_data = 12'hcff;
			{9'd86, 8'd122}: color_data = 12'h877;
			{9'd86, 8'd123}: color_data = 12'h002;
			{9'd86, 8'd124}: color_data = 12'h004;
			{9'd86, 8'd125}: color_data = 12'h004;
			{9'd86, 8'd126}: color_data = 12'h000;
			{9'd86, 8'd127}: color_data = 12'h068;
			{9'd86, 8'd128}: color_data = 12'h079;
			{9'd86, 8'd129}: color_data = 12'h000;
			{9'd86, 8'd170}: color_data = 12'h000;
			{9'd86, 8'd171}: color_data = 12'h068;
			{9'd86, 8'd172}: color_data = 12'h8ff;
			{9'd86, 8'd173}: color_data = 12'hcbb;
			{9'd86, 8'd174}: color_data = 12'h323;
			{9'd86, 8'd175}: color_data = 12'h003;
			{9'd86, 8'd176}: color_data = 12'h005;
			{9'd86, 8'd177}: color_data = 12'h002;
			{9'd86, 8'd178}: color_data = 12'h023;
			{9'd86, 8'd179}: color_data = 12'h09c;
			{9'd86, 8'd180}: color_data = 12'h023;
			{9'd86, 8'd222}: color_data = 12'h100;
			{9'd86, 8'd223}: color_data = 12'h800;
			{9'd86, 8'd224}: color_data = 12'h900;
			{9'd86, 8'd225}: color_data = 12'h800;
			{9'd86, 8'd226}: color_data = 12'h100;
			{9'd86, 8'd227}: color_data = 12'h510;
			{9'd86, 8'd228}: color_data = 12'h930;
			{9'd86, 8'd229}: color_data = 12'h610;
			{9'd86, 8'd230}: color_data = 12'h100;
			{9'd86, 8'd231}: color_data = 12'h300;
			{9'd86, 8'd232}: color_data = 12'h900;
			{9'd86, 8'd233}: color_data = 12'ha00;
			{9'd86, 8'd234}: color_data = 12'h600;
			{9'd86, 8'd235}: color_data = 12'h100;
			{9'd86, 8'd236}: color_data = 12'h820;
			{9'd86, 8'd237}: color_data = 12'h920;
			{9'd86, 8'd238}: color_data = 12'h500;
			{9'd86, 8'd239}: color_data = 12'h000;
			{9'd87, 8'd68}: color_data = 12'h057;
			{9'd87, 8'd69}: color_data = 12'h3bd;
			{9'd87, 8'd70}: color_data = 12'h555;
			{9'd87, 8'd71}: color_data = 12'h002;
			{9'd87, 8'd72}: color_data = 12'h005;
			{9'd87, 8'd73}: color_data = 12'h005;
			{9'd87, 8'd74}: color_data = 12'h004;
			{9'd87, 8'd75}: color_data = 12'h025;
			{9'd87, 8'd76}: color_data = 12'h09c;
			{9'd87, 8'd77}: color_data = 12'h034;
			{9'd87, 8'd119}: color_data = 12'h000;
			{9'd87, 8'd120}: color_data = 12'h1ac;
			{9'd87, 8'd121}: color_data = 12'h689;
			{9'd87, 8'd122}: color_data = 12'h212;
			{9'd87, 8'd123}: color_data = 12'h004;
			{9'd87, 8'd124}: color_data = 12'h005;
			{9'd87, 8'd125}: color_data = 12'h005;
			{9'd87, 8'd126}: color_data = 12'h003;
			{9'd87, 8'd127}: color_data = 12'h06a;
			{9'd87, 8'd128}: color_data = 12'h079;
			{9'd87, 8'd129}: color_data = 12'h000;
			{9'd87, 8'd170}: color_data = 12'h000;
			{9'd87, 8'd171}: color_data = 12'h079;
			{9'd87, 8'd172}: color_data = 12'h4bd;
			{9'd87, 8'd173}: color_data = 12'h444;
			{9'd87, 8'd174}: color_data = 12'h002;
			{9'd87, 8'd175}: color_data = 12'h005;
			{9'd87, 8'd176}: color_data = 12'h005;
			{9'd87, 8'd177}: color_data = 12'h004;
			{9'd87, 8'd178}: color_data = 12'h036;
			{9'd87, 8'd179}: color_data = 12'h09c;
			{9'd87, 8'd180}: color_data = 12'h023;
			{9'd87, 8'd222}: color_data = 12'h200;
			{9'd87, 8'd223}: color_data = 12'ha00;
			{9'd87, 8'd224}: color_data = 12'ha00;
			{9'd87, 8'd225}: color_data = 12'h800;
			{9'd87, 8'd226}: color_data = 12'h100;
			{9'd87, 8'd227}: color_data = 12'h100;
			{9'd87, 8'd228}: color_data = 12'h200;
			{9'd87, 8'd229}: color_data = 12'h200;
			{9'd87, 8'd230}: color_data = 12'h000;
			{9'd87, 8'd231}: color_data = 12'h500;
			{9'd87, 8'd232}: color_data = 12'hb00;
			{9'd87, 8'd233}: color_data = 12'ha00;
			{9'd87, 8'd234}: color_data = 12'h700;
			{9'd87, 8'd235}: color_data = 12'h000;
			{9'd87, 8'd236}: color_data = 12'h100;
			{9'd87, 8'd237}: color_data = 12'h200;
			{9'd87, 8'd238}: color_data = 12'h200;
			{9'd87, 8'd239}: color_data = 12'h100;
			{9'd88, 8'd68}: color_data = 12'h035;
			{9'd88, 8'd69}: color_data = 12'h047;
			{9'd88, 8'd70}: color_data = 12'h001;
			{9'd88, 8'd71}: color_data = 12'h004;
			{9'd88, 8'd72}: color_data = 12'h004;
			{9'd88, 8'd73}: color_data = 12'h004;
			{9'd88, 8'd74}: color_data = 12'h004;
			{9'd88, 8'd75}: color_data = 12'h015;
			{9'd88, 8'd76}: color_data = 12'h059;
			{9'd88, 8'd77}: color_data = 12'h023;
			{9'd88, 8'd119}: color_data = 12'h000;
			{9'd88, 8'd120}: color_data = 12'h058;
			{9'd88, 8'd121}: color_data = 12'h013;
			{9'd88, 8'd122}: color_data = 12'h002;
			{9'd88, 8'd123}: color_data = 12'h004;
			{9'd88, 8'd124}: color_data = 12'h004;
			{9'd88, 8'd125}: color_data = 12'h004;
			{9'd88, 8'd126}: color_data = 12'h004;
			{9'd88, 8'd127}: color_data = 12'h038;
			{9'd88, 8'd128}: color_data = 12'h046;
			{9'd88, 8'd129}: color_data = 12'h000;
			{9'd88, 8'd170}: color_data = 12'h000;
			{9'd88, 8'd171}: color_data = 12'h047;
			{9'd88, 8'd172}: color_data = 12'h036;
			{9'd88, 8'd173}: color_data = 12'h001;
			{9'd88, 8'd174}: color_data = 12'h004;
			{9'd88, 8'd175}: color_data = 12'h004;
			{9'd88, 8'd176}: color_data = 12'h004;
			{9'd88, 8'd177}: color_data = 12'h004;
			{9'd88, 8'd178}: color_data = 12'h016;
			{9'd88, 8'd179}: color_data = 12'h059;
			{9'd88, 8'd180}: color_data = 12'h012;
			{9'd88, 8'd222}: color_data = 12'h410;
			{9'd88, 8'd223}: color_data = 12'he40;
			{9'd88, 8'd224}: color_data = 12'hd20;
			{9'd88, 8'd225}: color_data = 12'h900;
			{9'd88, 8'd226}: color_data = 12'h200;
			{9'd88, 8'd227}: color_data = 12'h600;
			{9'd88, 8'd228}: color_data = 12'ha00;
			{9'd88, 8'd229}: color_data = 12'h900;
			{9'd88, 8'd230}: color_data = 12'h200;
			{9'd88, 8'd231}: color_data = 12'h820;
			{9'd88, 8'd232}: color_data = 12'hf30;
			{9'd88, 8'd233}: color_data = 12'hc00;
			{9'd88, 8'd234}: color_data = 12'h500;
			{9'd88, 8'd235}: color_data = 12'h200;
			{9'd88, 8'd236}: color_data = 12'h800;
			{9'd88, 8'd237}: color_data = 12'ha00;
			{9'd88, 8'd238}: color_data = 12'h700;
			{9'd88, 8'd239}: color_data = 12'h100;
			{9'd89, 8'd68}: color_data = 12'h013;
			{9'd89, 8'd69}: color_data = 12'h027;
			{9'd89, 8'd70}: color_data = 12'h016;
			{9'd89, 8'd71}: color_data = 12'h027;
			{9'd89, 8'd72}: color_data = 12'h027;
			{9'd89, 8'd73}: color_data = 12'h026;
			{9'd89, 8'd74}: color_data = 12'h027;
			{9'd89, 8'd75}: color_data = 12'h028;
			{9'd89, 8'd76}: color_data = 12'h027;
			{9'd89, 8'd77}: color_data = 12'h001;
			{9'd89, 8'd119}: color_data = 12'h000;
			{9'd89, 8'd120}: color_data = 12'h016;
			{9'd89, 8'd121}: color_data = 12'h017;
			{9'd89, 8'd122}: color_data = 12'h016;
			{9'd89, 8'd123}: color_data = 12'h027;
			{9'd89, 8'd124}: color_data = 12'h027;
			{9'd89, 8'd125}: color_data = 12'h027;
			{9'd89, 8'd126}: color_data = 12'h027;
			{9'd89, 8'd127}: color_data = 12'h028;
			{9'd89, 8'd128}: color_data = 12'h014;
			{9'd89, 8'd129}: color_data = 12'h000;
			{9'd89, 8'd170}: color_data = 12'h000;
			{9'd89, 8'd171}: color_data = 12'h014;
			{9'd89, 8'd172}: color_data = 12'h027;
			{9'd89, 8'd173}: color_data = 12'h016;
			{9'd89, 8'd174}: color_data = 12'h027;
			{9'd89, 8'd175}: color_data = 12'h027;
			{9'd89, 8'd176}: color_data = 12'h026;
			{9'd89, 8'd177}: color_data = 12'h027;
			{9'd89, 8'd178}: color_data = 12'h028;
			{9'd89, 8'd179}: color_data = 12'h026;
			{9'd89, 8'd180}: color_data = 12'h001;
			{9'd89, 8'd222}: color_data = 12'h300;
			{9'd89, 8'd223}: color_data = 12'hc30;
			{9'd89, 8'd224}: color_data = 12'hc30;
			{9'd89, 8'd225}: color_data = 12'h600;
			{9'd89, 8'd226}: color_data = 12'h100;
			{9'd89, 8'd227}: color_data = 12'h600;
			{9'd89, 8'd228}: color_data = 12'ha00;
			{9'd89, 8'd229}: color_data = 12'h900;
			{9'd89, 8'd230}: color_data = 12'h300;
			{9'd89, 8'd231}: color_data = 12'h620;
			{9'd89, 8'd232}: color_data = 12'hd40;
			{9'd89, 8'd233}: color_data = 12'ha20;
			{9'd89, 8'd234}: color_data = 12'h300;
			{9'd89, 8'd235}: color_data = 12'h200;
			{9'd89, 8'd236}: color_data = 12'h900;
			{9'd89, 8'd237}: color_data = 12'ha00;
			{9'd89, 8'd238}: color_data = 12'h700;
			{9'd89, 8'd239}: color_data = 12'h100;
			{9'd90, 8'd68}: color_data = 12'h035;
			{9'd90, 8'd69}: color_data = 12'h09e;
			{9'd90, 8'd70}: color_data = 12'h09e;
			{9'd90, 8'd71}: color_data = 12'h09e;
			{9'd90, 8'd72}: color_data = 12'h09e;
			{9'd90, 8'd73}: color_data = 12'h09e;
			{9'd90, 8'd74}: color_data = 12'h09e;
			{9'd90, 8'd75}: color_data = 12'h09e;
			{9'd90, 8'd76}: color_data = 12'h08c;
			{9'd90, 8'd77}: color_data = 12'h023;
			{9'd90, 8'd119}: color_data = 12'h000;
			{9'd90, 8'd120}: color_data = 12'h07b;
			{9'd90, 8'd121}: color_data = 12'h0ae;
			{9'd90, 8'd122}: color_data = 12'h09e;
			{9'd90, 8'd123}: color_data = 12'h09e;
			{9'd90, 8'd124}: color_data = 12'h09e;
			{9'd90, 8'd125}: color_data = 12'h09e;
			{9'd90, 8'd126}: color_data = 12'h09e;
			{9'd90, 8'd127}: color_data = 12'h09e;
			{9'd90, 8'd128}: color_data = 12'h057;
			{9'd90, 8'd129}: color_data = 12'h000;
			{9'd90, 8'd170}: color_data = 12'h000;
			{9'd90, 8'd171}: color_data = 12'h057;
			{9'd90, 8'd172}: color_data = 12'h0ae;
			{9'd90, 8'd173}: color_data = 12'h09e;
			{9'd90, 8'd174}: color_data = 12'h09e;
			{9'd90, 8'd175}: color_data = 12'h09e;
			{9'd90, 8'd176}: color_data = 12'h09e;
			{9'd90, 8'd177}: color_data = 12'h09e;
			{9'd90, 8'd178}: color_data = 12'h09e;
			{9'd90, 8'd179}: color_data = 12'h07b;
			{9'd90, 8'd180}: color_data = 12'h012;
			{9'd90, 8'd222}: color_data = 12'h000;
			{9'd90, 8'd223}: color_data = 12'h200;
			{9'd90, 8'd224}: color_data = 12'h300;
			{9'd90, 8'd225}: color_data = 12'h100;
			{9'd90, 8'd226}: color_data = 12'h000;
			{9'd90, 8'd227}: color_data = 12'h700;
			{9'd90, 8'd228}: color_data = 12'ha00;
			{9'd90, 8'd229}: color_data = 12'h900;
			{9'd90, 8'd230}: color_data = 12'h300;
			{9'd90, 8'd231}: color_data = 12'h100;
			{9'd90, 8'd232}: color_data = 12'h310;
			{9'd90, 8'd233}: color_data = 12'h200;
			{9'd90, 8'd234}: color_data = 12'h000;
			{9'd90, 8'd235}: color_data = 12'h300;
			{9'd90, 8'd236}: color_data = 12'h900;
			{9'd90, 8'd237}: color_data = 12'ha00;
			{9'd90, 8'd238}: color_data = 12'h700;
			{9'd90, 8'd239}: color_data = 12'h100;
			{9'd91, 8'd68}: color_data = 12'h057;
			{9'd91, 8'd69}: color_data = 12'h4ef;
			{9'd91, 8'd70}: color_data = 12'h7ef;
			{9'd91, 8'd71}: color_data = 12'h0cf;
			{9'd91, 8'd72}: color_data = 12'h0cf;
			{9'd91, 8'd73}: color_data = 12'h0df;
			{9'd91, 8'd74}: color_data = 12'h0bd;
			{9'd91, 8'd75}: color_data = 12'h068;
			{9'd91, 8'd76}: color_data = 12'h09c;
			{9'd91, 8'd77}: color_data = 12'h034;
			{9'd91, 8'd119}: color_data = 12'h000;
			{9'd91, 8'd120}: color_data = 12'h1ad;
			{9'd91, 8'd121}: color_data = 12'h8ff;
			{9'd91, 8'd122}: color_data = 12'h3df;
			{9'd91, 8'd123}: color_data = 12'h0cf;
			{9'd91, 8'd124}: color_data = 12'h0cf;
			{9'd91, 8'd125}: color_data = 12'h0cf;
			{9'd91, 8'd126}: color_data = 12'h079;
			{9'd91, 8'd127}: color_data = 12'h08b;
			{9'd91, 8'd128}: color_data = 12'h079;
			{9'd91, 8'd129}: color_data = 12'h000;
			{9'd91, 8'd170}: color_data = 12'h000;
			{9'd91, 8'd171}: color_data = 12'h069;
			{9'd91, 8'd172}: color_data = 12'h6ef;
			{9'd91, 8'd173}: color_data = 12'h6ef;
			{9'd91, 8'd174}: color_data = 12'h0cf;
			{9'd91, 8'd175}: color_data = 12'h0cf;
			{9'd91, 8'd176}: color_data = 12'h0df;
			{9'd91, 8'd177}: color_data = 12'h0ac;
			{9'd91, 8'd178}: color_data = 12'h079;
			{9'd91, 8'd179}: color_data = 12'h09c;
			{9'd91, 8'd180}: color_data = 12'h023;
			{9'd91, 8'd222}: color_data = 12'h100;
			{9'd91, 8'd223}: color_data = 12'h400;
			{9'd91, 8'd224}: color_data = 12'h500;
			{9'd91, 8'd225}: color_data = 12'h400;
			{9'd91, 8'd226}: color_data = 12'h200;
			{9'd91, 8'd227}: color_data = 12'ha20;
			{9'd91, 8'd228}: color_data = 12'hb10;
			{9'd91, 8'd229}: color_data = 12'h900;
			{9'd91, 8'd230}: color_data = 12'h300;
			{9'd91, 8'd231}: color_data = 12'h200;
			{9'd91, 8'd232}: color_data = 12'h500;
			{9'd91, 8'd233}: color_data = 12'h500;
			{9'd91, 8'd234}: color_data = 12'h200;
			{9'd91, 8'd235}: color_data = 12'h410;
			{9'd91, 8'd236}: color_data = 12'hc20;
			{9'd91, 8'd237}: color_data = 12'ha00;
			{9'd91, 8'd238}: color_data = 12'h700;
			{9'd91, 8'd239}: color_data = 12'h100;
			{9'd92, 8'd68}: color_data = 12'h047;
			{9'd92, 8'd69}: color_data = 12'h6df;
			{9'd92, 8'd70}: color_data = 12'heff;
			{9'd92, 8'd71}: color_data = 12'h6df;
			{9'd92, 8'd72}: color_data = 12'h0bf;
			{9'd92, 8'd73}: color_data = 12'h0be;
			{9'd92, 8'd74}: color_data = 12'h056;
			{9'd92, 8'd75}: color_data = 12'h012;
			{9'd92, 8'd76}: color_data = 12'h08b;
			{9'd92, 8'd77}: color_data = 12'h034;
			{9'd92, 8'd119}: color_data = 12'h000;
			{9'd92, 8'd120}: color_data = 12'h2ac;
			{9'd92, 8'd121}: color_data = 12'hdff;
			{9'd92, 8'd122}: color_data = 12'haef;
			{9'd92, 8'd123}: color_data = 12'h1bf;
			{9'd92, 8'd124}: color_data = 12'h0cf;
			{9'd92, 8'd125}: color_data = 12'h08b;
			{9'd92, 8'd126}: color_data = 12'h012;
			{9'd92, 8'd127}: color_data = 12'h068;
			{9'd92, 8'd128}: color_data = 12'h079;
			{9'd92, 8'd129}: color_data = 12'h000;
			{9'd92, 8'd170}: color_data = 12'h000;
			{9'd92, 8'd171}: color_data = 12'h068;
			{9'd92, 8'd172}: color_data = 12'h8ef;
			{9'd92, 8'd173}: color_data = 12'hdff;
			{9'd92, 8'd174}: color_data = 12'h4cf;
			{9'd92, 8'd175}: color_data = 12'h0bf;
			{9'd92, 8'd176}: color_data = 12'h0ae;
			{9'd92, 8'd177}: color_data = 12'h035;
			{9'd92, 8'd178}: color_data = 12'h023;
			{9'd92, 8'd179}: color_data = 12'h08c;
			{9'd92, 8'd180}: color_data = 12'h023;
			{9'd92, 8'd222}: color_data = 12'h200;
			{9'd92, 8'd223}: color_data = 12'h900;
			{9'd92, 8'd224}: color_data = 12'hb00;
			{9'd92, 8'd225}: color_data = 12'h800;
			{9'd92, 8'd226}: color_data = 12'h200;
			{9'd92, 8'd227}: color_data = 12'hb30;
			{9'd92, 8'd228}: color_data = 12'hc10;
			{9'd92, 8'd229}: color_data = 12'h800;
			{9'd92, 8'd230}: color_data = 12'h300;
			{9'd92, 8'd231}: color_data = 12'h400;
			{9'd92, 8'd232}: color_data = 12'ha00;
			{9'd92, 8'd233}: color_data = 12'ha00;
			{9'd92, 8'd234}: color_data = 12'h500;
			{9'd92, 8'd235}: color_data = 12'h510;
			{9'd92, 8'd236}: color_data = 12'hd30;
			{9'd92, 8'd237}: color_data = 12'ha00;
			{9'd92, 8'd238}: color_data = 12'h700;
			{9'd92, 8'd239}: color_data = 12'h100;
			{9'd93, 8'd68}: color_data = 12'h047;
			{9'd93, 8'd69}: color_data = 12'h6df;
			{9'd93, 8'd70}: color_data = 12'hfff;
			{9'd93, 8'd71}: color_data = 12'hdff;
			{9'd93, 8'd72}: color_data = 12'h5df;
			{9'd93, 8'd73}: color_data = 12'h068;
			{9'd93, 8'd74}: color_data = 12'h000;
			{9'd93, 8'd75}: color_data = 12'h012;
			{9'd93, 8'd76}: color_data = 12'h08c;
			{9'd93, 8'd77}: color_data = 12'h034;
			{9'd93, 8'd119}: color_data = 12'h000;
			{9'd93, 8'd120}: color_data = 12'h1ac;
			{9'd93, 8'd121}: color_data = 12'hdff;
			{9'd93, 8'd122}: color_data = 12'hfff;
			{9'd93, 8'd123}: color_data = 12'h9ef;
			{9'd93, 8'd124}: color_data = 12'h19c;
			{9'd93, 8'd125}: color_data = 12'h023;
			{9'd93, 8'd127}: color_data = 12'h068;
			{9'd93, 8'd128}: color_data = 12'h079;
			{9'd93, 8'd129}: color_data = 12'h000;
			{9'd93, 8'd170}: color_data = 12'h000;
			{9'd93, 8'd171}: color_data = 12'h068;
			{9'd93, 8'd172}: color_data = 12'h8ef;
			{9'd93, 8'd173}: color_data = 12'hfff;
			{9'd93, 8'd174}: color_data = 12'hcff;
			{9'd93, 8'd175}: color_data = 12'h4ce;
			{9'd93, 8'd176}: color_data = 12'h057;
			{9'd93, 8'd177}: color_data = 12'h000;
			{9'd93, 8'd178}: color_data = 12'h023;
			{9'd93, 8'd179}: color_data = 12'h08c;
			{9'd93, 8'd180}: color_data = 12'h023;
			{9'd93, 8'd222}: color_data = 12'h200;
			{9'd93, 8'd223}: color_data = 12'h900;
			{9'd93, 8'd224}: color_data = 12'ha00;
			{9'd93, 8'd225}: color_data = 12'h700;
			{9'd93, 8'd226}: color_data = 12'h200;
			{9'd93, 8'd227}: color_data = 12'hb30;
			{9'd93, 8'd228}: color_data = 12'he20;
			{9'd93, 8'd229}: color_data = 12'ha00;
			{9'd93, 8'd230}: color_data = 12'h300;
			{9'd93, 8'd231}: color_data = 12'h400;
			{9'd93, 8'd232}: color_data = 12'ha00;
			{9'd93, 8'd233}: color_data = 12'ha00;
			{9'd93, 8'd234}: color_data = 12'h400;
			{9'd93, 8'd235}: color_data = 12'h510;
			{9'd93, 8'd236}: color_data = 12'hf40;
			{9'd93, 8'd237}: color_data = 12'hd10;
			{9'd93, 8'd238}: color_data = 12'h800;
			{9'd93, 8'd239}: color_data = 12'h100;
			{9'd94, 8'd68}: color_data = 12'h047;
			{9'd94, 8'd69}: color_data = 12'h6df;
			{9'd94, 8'd70}: color_data = 12'hfff;
			{9'd94, 8'd71}: color_data = 12'hfff;
			{9'd94, 8'd72}: color_data = 12'h9aa;
			{9'd94, 8'd73}: color_data = 12'h011;
			{9'd94, 8'd75}: color_data = 12'h012;
			{9'd94, 8'd76}: color_data = 12'h08c;
			{9'd94, 8'd77}: color_data = 12'h034;
			{9'd94, 8'd119}: color_data = 12'h000;
			{9'd94, 8'd120}: color_data = 12'h1ac;
			{9'd94, 8'd121}: color_data = 12'hcff;
			{9'd94, 8'd122}: color_data = 12'hfff;
			{9'd94, 8'd123}: color_data = 12'hddd;
			{9'd94, 8'd124}: color_data = 12'h345;
			{9'd94, 8'd126}: color_data = 12'h000;
			{9'd94, 8'd127}: color_data = 12'h068;
			{9'd94, 8'd128}: color_data = 12'h079;
			{9'd94, 8'd129}: color_data = 12'h000;
			{9'd94, 8'd170}: color_data = 12'h000;
			{9'd94, 8'd171}: color_data = 12'h068;
			{9'd94, 8'd172}: color_data = 12'h7ef;
			{9'd94, 8'd173}: color_data = 12'hfff;
			{9'd94, 8'd174}: color_data = 12'hfff;
			{9'd94, 8'd175}: color_data = 12'h899;
			{9'd94, 8'd176}: color_data = 12'h001;
			{9'd94, 8'd178}: color_data = 12'h024;
			{9'd94, 8'd179}: color_data = 12'h08c;
			{9'd94, 8'd180}: color_data = 12'h023;
			{9'd94, 8'd222}: color_data = 12'h200;
			{9'd94, 8'd223}: color_data = 12'h800;
			{9'd94, 8'd224}: color_data = 12'ha00;
			{9'd94, 8'd225}: color_data = 12'h700;
			{9'd94, 8'd226}: color_data = 12'h200;
			{9'd94, 8'd227}: color_data = 12'h920;
			{9'd94, 8'd228}: color_data = 12'hd30;
			{9'd94, 8'd229}: color_data = 12'h910;
			{9'd94, 8'd230}: color_data = 12'h200;
			{9'd94, 8'd231}: color_data = 12'h400;
			{9'd94, 8'd232}: color_data = 12'h900;
			{9'd94, 8'd233}: color_data = 12'ha00;
			{9'd94, 8'd234}: color_data = 12'h400;
			{9'd94, 8'd235}: color_data = 12'h310;
			{9'd94, 8'd236}: color_data = 12'hc30;
			{9'd94, 8'd237}: color_data = 12'hc20;
			{9'd94, 8'd238}: color_data = 12'h600;
			{9'd94, 8'd239}: color_data = 12'h000;
			{9'd95, 8'd68}: color_data = 12'h047;
			{9'd95, 8'd69}: color_data = 12'h6df;
			{9'd95, 8'd70}: color_data = 12'hfff;
			{9'd95, 8'd71}: color_data = 12'hcbb;
			{9'd95, 8'd72}: color_data = 12'h323;
			{9'd95, 8'd73}: color_data = 12'h002;
			{9'd95, 8'd74}: color_data = 12'h000;
			{9'd95, 8'd75}: color_data = 12'h012;
			{9'd95, 8'd76}: color_data = 12'h08c;
			{9'd95, 8'd77}: color_data = 12'h034;
			{9'd95, 8'd119}: color_data = 12'h000;
			{9'd95, 8'd120}: color_data = 12'h1ac;
			{9'd95, 8'd121}: color_data = 12'hdff;
			{9'd95, 8'd122}: color_data = 12'hfee;
			{9'd95, 8'd123}: color_data = 12'h666;
			{9'd95, 8'd124}: color_data = 12'h002;
			{9'd95, 8'd125}: color_data = 12'h001;
			{9'd95, 8'd126}: color_data = 12'h000;
			{9'd95, 8'd127}: color_data = 12'h068;
			{9'd95, 8'd128}: color_data = 12'h079;
			{9'd95, 8'd129}: color_data = 12'h000;
			{9'd95, 8'd170}: color_data = 12'h000;
			{9'd95, 8'd171}: color_data = 12'h068;
			{9'd95, 8'd172}: color_data = 12'h8ef;
			{9'd95, 8'd173}: color_data = 12'hfff;
			{9'd95, 8'd174}: color_data = 12'haaa;
			{9'd95, 8'd175}: color_data = 12'h212;
			{9'd95, 8'd176}: color_data = 12'h002;
			{9'd95, 8'd178}: color_data = 12'h023;
			{9'd95, 8'd179}: color_data = 12'h08c;
			{9'd95, 8'd180}: color_data = 12'h023;
			{9'd95, 8'd222}: color_data = 12'h200;
			{9'd95, 8'd223}: color_data = 12'h900;
			{9'd95, 8'd224}: color_data = 12'ha00;
			{9'd95, 8'd225}: color_data = 12'h800;
			{9'd95, 8'd226}: color_data = 12'h100;
			{9'd95, 8'd227}: color_data = 12'h100;
			{9'd95, 8'd228}: color_data = 12'h310;
			{9'd95, 8'd229}: color_data = 12'h200;
			{9'd95, 8'd230}: color_data = 12'h000;
			{9'd95, 8'd231}: color_data = 12'h500;
			{9'd95, 8'd232}: color_data = 12'ha00;
			{9'd95, 8'd233}: color_data = 12'ha00;
			{9'd95, 8'd234}: color_data = 12'h500;
			{9'd95, 8'd235}: color_data = 12'h000;
			{9'd95, 8'd236}: color_data = 12'h200;
			{9'd95, 8'd237}: color_data = 12'h300;
			{9'd95, 8'd238}: color_data = 12'h100;
			{9'd95, 8'd239}: color_data = 12'h000;
			{9'd96, 8'd68}: color_data = 12'h047;
			{9'd96, 8'd69}: color_data = 12'h6ef;
			{9'd96, 8'd70}: color_data = 12'hddc;
			{9'd96, 8'd71}: color_data = 12'h434;
			{9'd96, 8'd72}: color_data = 12'h003;
			{9'd96, 8'd73}: color_data = 12'h005;
			{9'd96, 8'd74}: color_data = 12'h002;
			{9'd96, 8'd75}: color_data = 12'h012;
			{9'd96, 8'd76}: color_data = 12'h08c;
			{9'd96, 8'd77}: color_data = 12'h034;
			{9'd96, 8'd119}: color_data = 12'h000;
			{9'd96, 8'd120}: color_data = 12'h2ad;
			{9'd96, 8'd121}: color_data = 12'hcff;
			{9'd96, 8'd122}: color_data = 12'h877;
			{9'd96, 8'd123}: color_data = 12'h002;
			{9'd96, 8'd124}: color_data = 12'h004;
			{9'd96, 8'd125}: color_data = 12'h004;
			{9'd96, 8'd126}: color_data = 12'h000;
			{9'd96, 8'd127}: color_data = 12'h068;
			{9'd96, 8'd128}: color_data = 12'h079;
			{9'd96, 8'd129}: color_data = 12'h000;
			{9'd96, 8'd170}: color_data = 12'h000;
			{9'd96, 8'd171}: color_data = 12'h068;
			{9'd96, 8'd172}: color_data = 12'h8ff;
			{9'd96, 8'd173}: color_data = 12'hcbb;
			{9'd96, 8'd174}: color_data = 12'h223;
			{9'd96, 8'd175}: color_data = 12'h003;
			{9'd96, 8'd176}: color_data = 12'h005;
			{9'd96, 8'd177}: color_data = 12'h002;
			{9'd96, 8'd178}: color_data = 12'h023;
			{9'd96, 8'd179}: color_data = 12'h09c;
			{9'd96, 8'd180}: color_data = 12'h023;
			{9'd96, 8'd222}: color_data = 12'h300;
			{9'd96, 8'd223}: color_data = 12'hc20;
			{9'd96, 8'd224}: color_data = 12'ha00;
			{9'd96, 8'd225}: color_data = 12'h800;
			{9'd96, 8'd226}: color_data = 12'h100;
			{9'd96, 8'd227}: color_data = 12'h300;
			{9'd96, 8'd228}: color_data = 12'h500;
			{9'd96, 8'd229}: color_data = 12'h500;
			{9'd96, 8'd230}: color_data = 12'h100;
			{9'd96, 8'd231}: color_data = 12'h710;
			{9'd96, 8'd232}: color_data = 12'hc10;
			{9'd96, 8'd233}: color_data = 12'h900;
			{9'd96, 8'd234}: color_data = 12'h500;
			{9'd96, 8'd235}: color_data = 12'h100;
			{9'd96, 8'd236}: color_data = 12'h500;
			{9'd96, 8'd237}: color_data = 12'h500;
			{9'd96, 8'd238}: color_data = 12'h400;
			{9'd96, 8'd239}: color_data = 12'h000;
			{9'd97, 8'd68}: color_data = 12'h057;
			{9'd97, 8'd69}: color_data = 12'h3bd;
			{9'd97, 8'd70}: color_data = 12'h555;
			{9'd97, 8'd71}: color_data = 12'h002;
			{9'd97, 8'd72}: color_data = 12'h005;
			{9'd97, 8'd73}: color_data = 12'h005;
			{9'd97, 8'd74}: color_data = 12'h004;
			{9'd97, 8'd75}: color_data = 12'h025;
			{9'd97, 8'd76}: color_data = 12'h09c;
			{9'd97, 8'd77}: color_data = 12'h034;
			{9'd97, 8'd119}: color_data = 12'h000;
			{9'd97, 8'd120}: color_data = 12'h1ac;
			{9'd97, 8'd121}: color_data = 12'h699;
			{9'd97, 8'd122}: color_data = 12'h212;
			{9'd97, 8'd123}: color_data = 12'h004;
			{9'd97, 8'd124}: color_data = 12'h005;
			{9'd97, 8'd125}: color_data = 12'h005;
			{9'd97, 8'd126}: color_data = 12'h003;
			{9'd97, 8'd127}: color_data = 12'h06a;
			{9'd97, 8'd128}: color_data = 12'h079;
			{9'd97, 8'd129}: color_data = 12'h000;
			{9'd97, 8'd170}: color_data = 12'h000;
			{9'd97, 8'd171}: color_data = 12'h079;
			{9'd97, 8'd172}: color_data = 12'h4bd;
			{9'd97, 8'd173}: color_data = 12'h444;
			{9'd97, 8'd174}: color_data = 12'h002;
			{9'd97, 8'd175}: color_data = 12'h005;
			{9'd97, 8'd176}: color_data = 12'h005;
			{9'd97, 8'd177}: color_data = 12'h004;
			{9'd97, 8'd178}: color_data = 12'h036;
			{9'd97, 8'd179}: color_data = 12'h09c;
			{9'd97, 8'd180}: color_data = 12'h023;
			{9'd97, 8'd222}: color_data = 12'h410;
			{9'd97, 8'd223}: color_data = 12'hd30;
			{9'd97, 8'd224}: color_data = 12'hb00;
			{9'd97, 8'd225}: color_data = 12'h700;
			{9'd97, 8'd226}: color_data = 12'h200;
			{9'd97, 8'd227}: color_data = 12'h700;
			{9'd97, 8'd228}: color_data = 12'hb00;
			{9'd97, 8'd229}: color_data = 12'ha00;
			{9'd97, 8'd230}: color_data = 12'h300;
			{9'd97, 8'd231}: color_data = 12'h820;
			{9'd97, 8'd232}: color_data = 12'hd20;
			{9'd97, 8'd233}: color_data = 12'h900;
			{9'd97, 8'd234}: color_data = 12'h500;
			{9'd97, 8'd235}: color_data = 12'h300;
			{9'd97, 8'd236}: color_data = 12'h900;
			{9'd97, 8'd237}: color_data = 12'hb00;
			{9'd97, 8'd238}: color_data = 12'h800;
			{9'd97, 8'd239}: color_data = 12'h100;
			{9'd98, 8'd68}: color_data = 12'h036;
			{9'd98, 8'd69}: color_data = 12'h047;
			{9'd98, 8'd70}: color_data = 12'h001;
			{9'd98, 8'd71}: color_data = 12'h004;
			{9'd98, 8'd72}: color_data = 12'h004;
			{9'd98, 8'd73}: color_data = 12'h004;
			{9'd98, 8'd74}: color_data = 12'h004;
			{9'd98, 8'd75}: color_data = 12'h015;
			{9'd98, 8'd76}: color_data = 12'h059;
			{9'd98, 8'd77}: color_data = 12'h023;
			{9'd98, 8'd119}: color_data = 12'h000;
			{9'd98, 8'd120}: color_data = 12'h058;
			{9'd98, 8'd121}: color_data = 12'h013;
			{9'd98, 8'd122}: color_data = 12'h002;
			{9'd98, 8'd123}: color_data = 12'h004;
			{9'd98, 8'd124}: color_data = 12'h004;
			{9'd98, 8'd125}: color_data = 12'h004;
			{9'd98, 8'd126}: color_data = 12'h004;
			{9'd98, 8'd127}: color_data = 12'h039;
			{9'd98, 8'd128}: color_data = 12'h046;
			{9'd98, 8'd129}: color_data = 12'h000;
			{9'd98, 8'd170}: color_data = 12'h000;
			{9'd98, 8'd171}: color_data = 12'h047;
			{9'd98, 8'd172}: color_data = 12'h036;
			{9'd98, 8'd173}: color_data = 12'h001;
			{9'd98, 8'd174}: color_data = 12'h004;
			{9'd98, 8'd175}: color_data = 12'h004;
			{9'd98, 8'd176}: color_data = 12'h004;
			{9'd98, 8'd177}: color_data = 12'h004;
			{9'd98, 8'd178}: color_data = 12'h016;
			{9'd98, 8'd179}: color_data = 12'h059;
			{9'd98, 8'd180}: color_data = 12'h012;
			{9'd98, 8'd222}: color_data = 12'h410;
			{9'd98, 8'd223}: color_data = 12'he40;
			{9'd98, 8'd224}: color_data = 12'hd20;
			{9'd98, 8'd225}: color_data = 12'h800;
			{9'd98, 8'd226}: color_data = 12'h200;
			{9'd98, 8'd227}: color_data = 12'h600;
			{9'd98, 8'd228}: color_data = 12'ha00;
			{9'd98, 8'd229}: color_data = 12'h900;
			{9'd98, 8'd230}: color_data = 12'h300;
			{9'd98, 8'd231}: color_data = 12'h820;
			{9'd98, 8'd232}: color_data = 12'hf30;
			{9'd98, 8'd233}: color_data = 12'hc00;
			{9'd98, 8'd234}: color_data = 12'h500;
			{9'd98, 8'd235}: color_data = 12'h200;
			{9'd98, 8'd236}: color_data = 12'h900;
			{9'd98, 8'd237}: color_data = 12'ha00;
			{9'd98, 8'd238}: color_data = 12'h700;
			{9'd98, 8'd239}: color_data = 12'h100;
			{9'd99, 8'd68}: color_data = 12'h013;
			{9'd99, 8'd69}: color_data = 12'h027;
			{9'd99, 8'd70}: color_data = 12'h016;
			{9'd99, 8'd71}: color_data = 12'h027;
			{9'd99, 8'd72}: color_data = 12'h027;
			{9'd99, 8'd73}: color_data = 12'h017;
			{9'd99, 8'd74}: color_data = 12'h027;
			{9'd99, 8'd75}: color_data = 12'h028;
			{9'd99, 8'd76}: color_data = 12'h027;
			{9'd99, 8'd77}: color_data = 12'h001;
			{9'd99, 8'd119}: color_data = 12'h000;
			{9'd99, 8'd120}: color_data = 12'h016;
			{9'd99, 8'd121}: color_data = 12'h017;
			{9'd99, 8'd122}: color_data = 12'h016;
			{9'd99, 8'd123}: color_data = 12'h027;
			{9'd99, 8'd124}: color_data = 12'h027;
			{9'd99, 8'd125}: color_data = 12'h017;
			{9'd99, 8'd126}: color_data = 12'h027;
			{9'd99, 8'd127}: color_data = 12'h028;
			{9'd99, 8'd128}: color_data = 12'h014;
			{9'd99, 8'd129}: color_data = 12'h000;
			{9'd99, 8'd170}: color_data = 12'h000;
			{9'd99, 8'd171}: color_data = 12'h014;
			{9'd99, 8'd172}: color_data = 12'h027;
			{9'd99, 8'd173}: color_data = 12'h016;
			{9'd99, 8'd174}: color_data = 12'h027;
			{9'd99, 8'd175}: color_data = 12'h027;
			{9'd99, 8'd176}: color_data = 12'h017;
			{9'd99, 8'd177}: color_data = 12'h027;
			{9'd99, 8'd178}: color_data = 12'h028;
			{9'd99, 8'd179}: color_data = 12'h026;
			{9'd99, 8'd180}: color_data = 12'h001;
			{9'd99, 8'd222}: color_data = 12'h300;
			{9'd99, 8'd223}: color_data = 12'hc30;
			{9'd99, 8'd224}: color_data = 12'hc30;
			{9'd99, 8'd225}: color_data = 12'h700;
			{9'd99, 8'd226}: color_data = 12'h100;
			{9'd99, 8'd227}: color_data = 12'h600;
			{9'd99, 8'd228}: color_data = 12'ha00;
			{9'd99, 8'd229}: color_data = 12'h900;
			{9'd99, 8'd230}: color_data = 12'h300;
			{9'd99, 8'd231}: color_data = 12'h620;
			{9'd99, 8'd232}: color_data = 12'hd40;
			{9'd99, 8'd233}: color_data = 12'ha20;
			{9'd99, 8'd234}: color_data = 12'h300;
			{9'd99, 8'd235}: color_data = 12'h200;
			{9'd99, 8'd236}: color_data = 12'h900;
			{9'd99, 8'd237}: color_data = 12'ha00;
			{9'd99, 8'd238}: color_data = 12'h700;
			{9'd99, 8'd239}: color_data = 12'h100;
			{9'd100, 8'd68}: color_data = 12'h035;
			{9'd100, 8'd69}: color_data = 12'h09e;
			{9'd100, 8'd70}: color_data = 12'h09e;
			{9'd100, 8'd71}: color_data = 12'h09e;
			{9'd100, 8'd72}: color_data = 12'h09e;
			{9'd100, 8'd73}: color_data = 12'h09e;
			{9'd100, 8'd74}: color_data = 12'h09e;
			{9'd100, 8'd75}: color_data = 12'h09e;
			{9'd100, 8'd76}: color_data = 12'h08c;
			{9'd100, 8'd77}: color_data = 12'h023;
			{9'd100, 8'd119}: color_data = 12'h000;
			{9'd100, 8'd120}: color_data = 12'h07b;
			{9'd100, 8'd121}: color_data = 12'h0ae;
			{9'd100, 8'd122}: color_data = 12'h09e;
			{9'd100, 8'd123}: color_data = 12'h09e;
			{9'd100, 8'd124}: color_data = 12'h09e;
			{9'd100, 8'd125}: color_data = 12'h09e;
			{9'd100, 8'd126}: color_data = 12'h09e;
			{9'd100, 8'd127}: color_data = 12'h09e;
			{9'd100, 8'd128}: color_data = 12'h057;
			{9'd100, 8'd129}: color_data = 12'h000;
			{9'd100, 8'd170}: color_data = 12'h000;
			{9'd100, 8'd171}: color_data = 12'h057;
			{9'd100, 8'd172}: color_data = 12'h0ae;
			{9'd100, 8'd173}: color_data = 12'h09e;
			{9'd100, 8'd174}: color_data = 12'h09e;
			{9'd100, 8'd175}: color_data = 12'h09e;
			{9'd100, 8'd176}: color_data = 12'h09e;
			{9'd100, 8'd177}: color_data = 12'h09e;
			{9'd100, 8'd178}: color_data = 12'h09e;
			{9'd100, 8'd179}: color_data = 12'h07b;
			{9'd100, 8'd180}: color_data = 12'h012;
			{9'd100, 8'd222}: color_data = 12'h000;
			{9'd100, 8'd223}: color_data = 12'h200;
			{9'd100, 8'd224}: color_data = 12'h300;
			{9'd100, 8'd225}: color_data = 12'h100;
			{9'd100, 8'd226}: color_data = 12'h000;
			{9'd100, 8'd227}: color_data = 12'h700;
			{9'd100, 8'd228}: color_data = 12'ha00;
			{9'd100, 8'd229}: color_data = 12'h900;
			{9'd100, 8'd230}: color_data = 12'h300;
			{9'd100, 8'd231}: color_data = 12'h100;
			{9'd100, 8'd232}: color_data = 12'h310;
			{9'd100, 8'd233}: color_data = 12'h200;
			{9'd100, 8'd234}: color_data = 12'h000;
			{9'd100, 8'd235}: color_data = 12'h300;
			{9'd100, 8'd236}: color_data = 12'h900;
			{9'd100, 8'd237}: color_data = 12'ha00;
			{9'd100, 8'd238}: color_data = 12'h700;
			{9'd100, 8'd239}: color_data = 12'h100;
			{9'd101, 8'd68}: color_data = 12'h057;
			{9'd101, 8'd69}: color_data = 12'h4ef;
			{9'd101, 8'd70}: color_data = 12'h7ef;
			{9'd101, 8'd71}: color_data = 12'h0cf;
			{9'd101, 8'd72}: color_data = 12'h0cf;
			{9'd101, 8'd73}: color_data = 12'h0df;
			{9'd101, 8'd74}: color_data = 12'h0bd;
			{9'd101, 8'd75}: color_data = 12'h068;
			{9'd101, 8'd76}: color_data = 12'h09c;
			{9'd101, 8'd77}: color_data = 12'h034;
			{9'd101, 8'd119}: color_data = 12'h000;
			{9'd101, 8'd120}: color_data = 12'h1ad;
			{9'd101, 8'd121}: color_data = 12'h8ff;
			{9'd101, 8'd122}: color_data = 12'h3df;
			{9'd101, 8'd123}: color_data = 12'h0cf;
			{9'd101, 8'd124}: color_data = 12'h0cf;
			{9'd101, 8'd125}: color_data = 12'h0cf;
			{9'd101, 8'd126}: color_data = 12'h07a;
			{9'd101, 8'd127}: color_data = 12'h08b;
			{9'd101, 8'd128}: color_data = 12'h079;
			{9'd101, 8'd129}: color_data = 12'h000;
			{9'd101, 8'd170}: color_data = 12'h000;
			{9'd101, 8'd171}: color_data = 12'h069;
			{9'd101, 8'd172}: color_data = 12'h6ef;
			{9'd101, 8'd173}: color_data = 12'h6ef;
			{9'd101, 8'd174}: color_data = 12'h0cf;
			{9'd101, 8'd175}: color_data = 12'h0cf;
			{9'd101, 8'd176}: color_data = 12'h0df;
			{9'd101, 8'd177}: color_data = 12'h0ad;
			{9'd101, 8'd178}: color_data = 12'h079;
			{9'd101, 8'd179}: color_data = 12'h09c;
			{9'd101, 8'd180}: color_data = 12'h023;
			{9'd101, 8'd222}: color_data = 12'h100;
			{9'd101, 8'd223}: color_data = 12'h400;
			{9'd101, 8'd224}: color_data = 12'h500;
			{9'd101, 8'd225}: color_data = 12'h400;
			{9'd101, 8'd226}: color_data = 12'h200;
			{9'd101, 8'd227}: color_data = 12'ha20;
			{9'd101, 8'd228}: color_data = 12'hb10;
			{9'd101, 8'd229}: color_data = 12'h900;
			{9'd101, 8'd230}: color_data = 12'h300;
			{9'd101, 8'd231}: color_data = 12'h200;
			{9'd101, 8'd232}: color_data = 12'h500;
			{9'd101, 8'd233}: color_data = 12'h500;
			{9'd101, 8'd234}: color_data = 12'h200;
			{9'd101, 8'd235}: color_data = 12'h410;
			{9'd101, 8'd236}: color_data = 12'hc20;
			{9'd101, 8'd237}: color_data = 12'ha00;
			{9'd101, 8'd238}: color_data = 12'h700;
			{9'd101, 8'd239}: color_data = 12'h100;
			{9'd102, 8'd68}: color_data = 12'h047;
			{9'd102, 8'd69}: color_data = 12'h6df;
			{9'd102, 8'd70}: color_data = 12'heff;
			{9'd102, 8'd71}: color_data = 12'h6df;
			{9'd102, 8'd72}: color_data = 12'h0bf;
			{9'd102, 8'd73}: color_data = 12'h0bf;
			{9'd102, 8'd74}: color_data = 12'h056;
			{9'd102, 8'd75}: color_data = 12'h012;
			{9'd102, 8'd76}: color_data = 12'h08b;
			{9'd102, 8'd77}: color_data = 12'h034;
			{9'd102, 8'd119}: color_data = 12'h000;
			{9'd102, 8'd120}: color_data = 12'h2ac;
			{9'd102, 8'd121}: color_data = 12'hdff;
			{9'd102, 8'd122}: color_data = 12'haef;
			{9'd102, 8'd123}: color_data = 12'h1bf;
			{9'd102, 8'd124}: color_data = 12'h0cf;
			{9'd102, 8'd125}: color_data = 12'h08b;
			{9'd102, 8'd126}: color_data = 12'h012;
			{9'd102, 8'd127}: color_data = 12'h068;
			{9'd102, 8'd128}: color_data = 12'h079;
			{9'd102, 8'd129}: color_data = 12'h000;
			{9'd102, 8'd170}: color_data = 12'h000;
			{9'd102, 8'd171}: color_data = 12'h068;
			{9'd102, 8'd172}: color_data = 12'h8ef;
			{9'd102, 8'd173}: color_data = 12'hdff;
			{9'd102, 8'd174}: color_data = 12'h4cf;
			{9'd102, 8'd175}: color_data = 12'h0bf;
			{9'd102, 8'd176}: color_data = 12'h0ae;
			{9'd102, 8'd177}: color_data = 12'h035;
			{9'd102, 8'd178}: color_data = 12'h023;
			{9'd102, 8'd179}: color_data = 12'h08c;
			{9'd102, 8'd180}: color_data = 12'h023;
			{9'd102, 8'd222}: color_data = 12'h200;
			{9'd102, 8'd223}: color_data = 12'h900;
			{9'd102, 8'd224}: color_data = 12'hb00;
			{9'd102, 8'd225}: color_data = 12'h800;
			{9'd102, 8'd226}: color_data = 12'h200;
			{9'd102, 8'd227}: color_data = 12'hb30;
			{9'd102, 8'd228}: color_data = 12'hc10;
			{9'd102, 8'd229}: color_data = 12'h800;
			{9'd102, 8'd230}: color_data = 12'h300;
			{9'd102, 8'd231}: color_data = 12'h500;
			{9'd102, 8'd232}: color_data = 12'ha00;
			{9'd102, 8'd233}: color_data = 12'ha00;
			{9'd102, 8'd234}: color_data = 12'h500;
			{9'd102, 8'd235}: color_data = 12'h510;
			{9'd102, 8'd236}: color_data = 12'hd30;
			{9'd102, 8'd237}: color_data = 12'ha00;
			{9'd102, 8'd238}: color_data = 12'h700;
			{9'd102, 8'd239}: color_data = 12'h100;
			{9'd103, 8'd68}: color_data = 12'h047;
			{9'd103, 8'd69}: color_data = 12'h6df;
			{9'd103, 8'd70}: color_data = 12'hfff;
			{9'd103, 8'd71}: color_data = 12'hdff;
			{9'd103, 8'd72}: color_data = 12'h5df;
			{9'd103, 8'd73}: color_data = 12'h068;
			{9'd103, 8'd74}: color_data = 12'h000;
			{9'd103, 8'd75}: color_data = 12'h012;
			{9'd103, 8'd76}: color_data = 12'h08c;
			{9'd103, 8'd77}: color_data = 12'h034;
			{9'd103, 8'd119}: color_data = 12'h000;
			{9'd103, 8'd120}: color_data = 12'h1ac;
			{9'd103, 8'd121}: color_data = 12'hdff;
			{9'd103, 8'd122}: color_data = 12'hfff;
			{9'd103, 8'd123}: color_data = 12'h8ef;
			{9'd103, 8'd124}: color_data = 12'h19c;
			{9'd103, 8'd125}: color_data = 12'h023;
			{9'd103, 8'd127}: color_data = 12'h068;
			{9'd103, 8'd128}: color_data = 12'h079;
			{9'd103, 8'd129}: color_data = 12'h000;
			{9'd103, 8'd170}: color_data = 12'h000;
			{9'd103, 8'd171}: color_data = 12'h068;
			{9'd103, 8'd172}: color_data = 12'h8ef;
			{9'd103, 8'd173}: color_data = 12'hfff;
			{9'd103, 8'd174}: color_data = 12'hcff;
			{9'd103, 8'd175}: color_data = 12'h4ce;
			{9'd103, 8'd176}: color_data = 12'h057;
			{9'd103, 8'd177}: color_data = 12'h000;
			{9'd103, 8'd178}: color_data = 12'h023;
			{9'd103, 8'd179}: color_data = 12'h08c;
			{9'd103, 8'd180}: color_data = 12'h023;
			{9'd103, 8'd222}: color_data = 12'h200;
			{9'd103, 8'd223}: color_data = 12'h900;
			{9'd103, 8'd224}: color_data = 12'ha00;
			{9'd103, 8'd225}: color_data = 12'h700;
			{9'd103, 8'd226}: color_data = 12'h200;
			{9'd103, 8'd227}: color_data = 12'hb30;
			{9'd103, 8'd228}: color_data = 12'he20;
			{9'd103, 8'd229}: color_data = 12'ha00;
			{9'd103, 8'd230}: color_data = 12'h300;
			{9'd103, 8'd231}: color_data = 12'h400;
			{9'd103, 8'd232}: color_data = 12'ha00;
			{9'd103, 8'd233}: color_data = 12'ha00;
			{9'd103, 8'd234}: color_data = 12'h400;
			{9'd103, 8'd235}: color_data = 12'h510;
			{9'd103, 8'd236}: color_data = 12'hf40;
			{9'd103, 8'd237}: color_data = 12'hd10;
			{9'd103, 8'd238}: color_data = 12'h800;
			{9'd103, 8'd239}: color_data = 12'h100;
			{9'd104, 8'd68}: color_data = 12'h047;
			{9'd104, 8'd69}: color_data = 12'h6df;
			{9'd104, 8'd70}: color_data = 12'hfff;
			{9'd104, 8'd71}: color_data = 12'hfff;
			{9'd104, 8'd72}: color_data = 12'h9aa;
			{9'd104, 8'd73}: color_data = 12'h011;
			{9'd104, 8'd75}: color_data = 12'h012;
			{9'd104, 8'd76}: color_data = 12'h08c;
			{9'd104, 8'd77}: color_data = 12'h034;
			{9'd104, 8'd119}: color_data = 12'h000;
			{9'd104, 8'd120}: color_data = 12'h1ac;
			{9'd104, 8'd121}: color_data = 12'hcff;
			{9'd104, 8'd122}: color_data = 12'hfff;
			{9'd104, 8'd123}: color_data = 12'hddd;
			{9'd104, 8'd124}: color_data = 12'h345;
			{9'd104, 8'd126}: color_data = 12'h000;
			{9'd104, 8'd127}: color_data = 12'h068;
			{9'd104, 8'd128}: color_data = 12'h079;
			{9'd104, 8'd129}: color_data = 12'h000;
			{9'd104, 8'd170}: color_data = 12'h000;
			{9'd104, 8'd171}: color_data = 12'h068;
			{9'd104, 8'd172}: color_data = 12'h7ef;
			{9'd104, 8'd173}: color_data = 12'hfff;
			{9'd104, 8'd174}: color_data = 12'hfff;
			{9'd104, 8'd175}: color_data = 12'h899;
			{9'd104, 8'd176}: color_data = 12'h001;
			{9'd104, 8'd178}: color_data = 12'h024;
			{9'd104, 8'd179}: color_data = 12'h08c;
			{9'd104, 8'd180}: color_data = 12'h023;
			{9'd104, 8'd222}: color_data = 12'h200;
			{9'd104, 8'd223}: color_data = 12'h800;
			{9'd104, 8'd224}: color_data = 12'ha00;
			{9'd104, 8'd225}: color_data = 12'h700;
			{9'd104, 8'd226}: color_data = 12'h200;
			{9'd104, 8'd227}: color_data = 12'h920;
			{9'd104, 8'd228}: color_data = 12'hd30;
			{9'd104, 8'd229}: color_data = 12'h910;
			{9'd104, 8'd230}: color_data = 12'h200;
			{9'd104, 8'd231}: color_data = 12'h400;
			{9'd104, 8'd232}: color_data = 12'h900;
			{9'd104, 8'd233}: color_data = 12'ha00;
			{9'd104, 8'd234}: color_data = 12'h400;
			{9'd104, 8'd235}: color_data = 12'h310;
			{9'd104, 8'd236}: color_data = 12'hc30;
			{9'd104, 8'd237}: color_data = 12'hc20;
			{9'd104, 8'd238}: color_data = 12'h600;
			{9'd104, 8'd239}: color_data = 12'h000;
			{9'd105, 8'd68}: color_data = 12'h047;
			{9'd105, 8'd69}: color_data = 12'h6df;
			{9'd105, 8'd70}: color_data = 12'hfff;
			{9'd105, 8'd71}: color_data = 12'hcbb;
			{9'd105, 8'd72}: color_data = 12'h323;
			{9'd105, 8'd73}: color_data = 12'h002;
			{9'd105, 8'd74}: color_data = 12'h000;
			{9'd105, 8'd75}: color_data = 12'h012;
			{9'd105, 8'd76}: color_data = 12'h08c;
			{9'd105, 8'd77}: color_data = 12'h034;
			{9'd105, 8'd119}: color_data = 12'h000;
			{9'd105, 8'd120}: color_data = 12'h1ac;
			{9'd105, 8'd121}: color_data = 12'hdff;
			{9'd105, 8'd122}: color_data = 12'hfee;
			{9'd105, 8'd123}: color_data = 12'h666;
			{9'd105, 8'd124}: color_data = 12'h002;
			{9'd105, 8'd125}: color_data = 12'h001;
			{9'd105, 8'd126}: color_data = 12'h000;
			{9'd105, 8'd127}: color_data = 12'h068;
			{9'd105, 8'd128}: color_data = 12'h079;
			{9'd105, 8'd129}: color_data = 12'h000;
			{9'd105, 8'd170}: color_data = 12'h000;
			{9'd105, 8'd171}: color_data = 12'h068;
			{9'd105, 8'd172}: color_data = 12'h8ef;
			{9'd105, 8'd173}: color_data = 12'hfff;
			{9'd105, 8'd174}: color_data = 12'haaa;
			{9'd105, 8'd175}: color_data = 12'h213;
			{9'd105, 8'd176}: color_data = 12'h002;
			{9'd105, 8'd178}: color_data = 12'h023;
			{9'd105, 8'd179}: color_data = 12'h08c;
			{9'd105, 8'd180}: color_data = 12'h023;
			{9'd105, 8'd222}: color_data = 12'h200;
			{9'd105, 8'd223}: color_data = 12'h900;
			{9'd105, 8'd224}: color_data = 12'ha00;
			{9'd105, 8'd225}: color_data = 12'h800;
			{9'd105, 8'd226}: color_data = 12'h100;
			{9'd105, 8'd227}: color_data = 12'h100;
			{9'd105, 8'd228}: color_data = 12'h310;
			{9'd105, 8'd229}: color_data = 12'h200;
			{9'd105, 8'd230}: color_data = 12'h000;
			{9'd105, 8'd231}: color_data = 12'h500;
			{9'd105, 8'd232}: color_data = 12'ha00;
			{9'd105, 8'd233}: color_data = 12'ha00;
			{9'd105, 8'd234}: color_data = 12'h500;
			{9'd105, 8'd235}: color_data = 12'h000;
			{9'd105, 8'd236}: color_data = 12'h200;
			{9'd105, 8'd237}: color_data = 12'h300;
			{9'd105, 8'd238}: color_data = 12'h100;
			{9'd105, 8'd239}: color_data = 12'h000;
			{9'd106, 8'd68}: color_data = 12'h047;
			{9'd106, 8'd69}: color_data = 12'h6ef;
			{9'd106, 8'd70}: color_data = 12'hdcc;
			{9'd106, 8'd71}: color_data = 12'h434;
			{9'd106, 8'd72}: color_data = 12'h003;
			{9'd106, 8'd73}: color_data = 12'h005;
			{9'd106, 8'd74}: color_data = 12'h002;
			{9'd106, 8'd75}: color_data = 12'h012;
			{9'd106, 8'd76}: color_data = 12'h08c;
			{9'd106, 8'd77}: color_data = 12'h034;
			{9'd106, 8'd119}: color_data = 12'h000;
			{9'd106, 8'd120}: color_data = 12'h2ad;
			{9'd106, 8'd121}: color_data = 12'hcff;
			{9'd106, 8'd122}: color_data = 12'h877;
			{9'd106, 8'd123}: color_data = 12'h002;
			{9'd106, 8'd124}: color_data = 12'h004;
			{9'd106, 8'd125}: color_data = 12'h004;
			{9'd106, 8'd126}: color_data = 12'h000;
			{9'd106, 8'd127}: color_data = 12'h068;
			{9'd106, 8'd128}: color_data = 12'h079;
			{9'd106, 8'd129}: color_data = 12'h000;
			{9'd106, 8'd170}: color_data = 12'h000;
			{9'd106, 8'd171}: color_data = 12'h068;
			{9'd106, 8'd172}: color_data = 12'h8ff;
			{9'd106, 8'd173}: color_data = 12'hcbb;
			{9'd106, 8'd174}: color_data = 12'h323;
			{9'd106, 8'd175}: color_data = 12'h003;
			{9'd106, 8'd176}: color_data = 12'h005;
			{9'd106, 8'd177}: color_data = 12'h002;
			{9'd106, 8'd178}: color_data = 12'h023;
			{9'd106, 8'd179}: color_data = 12'h09c;
			{9'd106, 8'd180}: color_data = 12'h023;
			{9'd106, 8'd222}: color_data = 12'h300;
			{9'd106, 8'd223}: color_data = 12'hc20;
			{9'd106, 8'd224}: color_data = 12'ha00;
			{9'd106, 8'd225}: color_data = 12'h800;
			{9'd106, 8'd226}: color_data = 12'h100;
			{9'd106, 8'd227}: color_data = 12'h300;
			{9'd106, 8'd228}: color_data = 12'h500;
			{9'd106, 8'd229}: color_data = 12'h500;
			{9'd106, 8'd230}: color_data = 12'h100;
			{9'd106, 8'd231}: color_data = 12'h710;
			{9'd106, 8'd232}: color_data = 12'hc10;
			{9'd106, 8'd233}: color_data = 12'h900;
			{9'd106, 8'd234}: color_data = 12'h500;
			{9'd106, 8'd235}: color_data = 12'h100;
			{9'd106, 8'd236}: color_data = 12'h500;
			{9'd106, 8'd237}: color_data = 12'h600;
			{9'd106, 8'd238}: color_data = 12'h400;
			{9'd106, 8'd239}: color_data = 12'h000;
			{9'd107, 8'd68}: color_data = 12'h057;
			{9'd107, 8'd69}: color_data = 12'h3bd;
			{9'd107, 8'd70}: color_data = 12'h555;
			{9'd107, 8'd71}: color_data = 12'h002;
			{9'd107, 8'd72}: color_data = 12'h005;
			{9'd107, 8'd73}: color_data = 12'h005;
			{9'd107, 8'd74}: color_data = 12'h004;
			{9'd107, 8'd75}: color_data = 12'h025;
			{9'd107, 8'd76}: color_data = 12'h09c;
			{9'd107, 8'd77}: color_data = 12'h034;
			{9'd107, 8'd119}: color_data = 12'h000;
			{9'd107, 8'd120}: color_data = 12'h1ac;
			{9'd107, 8'd121}: color_data = 12'h689;
			{9'd107, 8'd122}: color_data = 12'h212;
			{9'd107, 8'd123}: color_data = 12'h004;
			{9'd107, 8'd124}: color_data = 12'h005;
			{9'd107, 8'd125}: color_data = 12'h005;
			{9'd107, 8'd126}: color_data = 12'h003;
			{9'd107, 8'd127}: color_data = 12'h06a;
			{9'd107, 8'd128}: color_data = 12'h079;
			{9'd107, 8'd129}: color_data = 12'h000;
			{9'd107, 8'd170}: color_data = 12'h000;
			{9'd107, 8'd171}: color_data = 12'h079;
			{9'd107, 8'd172}: color_data = 12'h4bd;
			{9'd107, 8'd173}: color_data = 12'h444;
			{9'd107, 8'd174}: color_data = 12'h002;
			{9'd107, 8'd175}: color_data = 12'h005;
			{9'd107, 8'd176}: color_data = 12'h005;
			{9'd107, 8'd177}: color_data = 12'h004;
			{9'd107, 8'd178}: color_data = 12'h036;
			{9'd107, 8'd179}: color_data = 12'h09c;
			{9'd107, 8'd180}: color_data = 12'h023;
			{9'd107, 8'd222}: color_data = 12'h410;
			{9'd107, 8'd223}: color_data = 12'hd30;
			{9'd107, 8'd224}: color_data = 12'hb00;
			{9'd107, 8'd225}: color_data = 12'h700;
			{9'd107, 8'd226}: color_data = 12'h200;
			{9'd107, 8'd227}: color_data = 12'h700;
			{9'd107, 8'd228}: color_data = 12'hb00;
			{9'd107, 8'd229}: color_data = 12'ha00;
			{9'd107, 8'd230}: color_data = 12'h300;
			{9'd107, 8'd231}: color_data = 12'h820;
			{9'd107, 8'd232}: color_data = 12'hd20;
			{9'd107, 8'd233}: color_data = 12'h900;
			{9'd107, 8'd234}: color_data = 12'h500;
			{9'd107, 8'd235}: color_data = 12'h300;
			{9'd107, 8'd236}: color_data = 12'h900;
			{9'd107, 8'd237}: color_data = 12'hb00;
			{9'd107, 8'd238}: color_data = 12'h800;
			{9'd107, 8'd239}: color_data = 12'h100;
			{9'd108, 8'd68}: color_data = 12'h035;
			{9'd108, 8'd69}: color_data = 12'h047;
			{9'd108, 8'd70}: color_data = 12'h001;
			{9'd108, 8'd71}: color_data = 12'h004;
			{9'd108, 8'd72}: color_data = 12'h004;
			{9'd108, 8'd73}: color_data = 12'h004;
			{9'd108, 8'd74}: color_data = 12'h004;
			{9'd108, 8'd75}: color_data = 12'h015;
			{9'd108, 8'd76}: color_data = 12'h059;
			{9'd108, 8'd77}: color_data = 12'h023;
			{9'd108, 8'd119}: color_data = 12'h000;
			{9'd108, 8'd120}: color_data = 12'h058;
			{9'd108, 8'd121}: color_data = 12'h013;
			{9'd108, 8'd122}: color_data = 12'h002;
			{9'd108, 8'd123}: color_data = 12'h004;
			{9'd108, 8'd124}: color_data = 12'h004;
			{9'd108, 8'd125}: color_data = 12'h004;
			{9'd108, 8'd126}: color_data = 12'h004;
			{9'd108, 8'd127}: color_data = 12'h038;
			{9'd108, 8'd128}: color_data = 12'h046;
			{9'd108, 8'd129}: color_data = 12'h000;
			{9'd108, 8'd170}: color_data = 12'h000;
			{9'd108, 8'd171}: color_data = 12'h047;
			{9'd108, 8'd172}: color_data = 12'h047;
			{9'd108, 8'd173}: color_data = 12'h002;
			{9'd108, 8'd174}: color_data = 12'h005;
			{9'd108, 8'd175}: color_data = 12'h005;
			{9'd108, 8'd176}: color_data = 12'h005;
			{9'd108, 8'd177}: color_data = 12'h005;
			{9'd108, 8'd178}: color_data = 12'h017;
			{9'd108, 8'd179}: color_data = 12'h06a;
			{9'd108, 8'd180}: color_data = 12'h012;
			{9'd108, 8'd222}: color_data = 12'h410;
			{9'd108, 8'd223}: color_data = 12'he40;
			{9'd108, 8'd224}: color_data = 12'hd20;
			{9'd108, 8'd225}: color_data = 12'h800;
			{9'd108, 8'd226}: color_data = 12'h200;
			{9'd108, 8'd227}: color_data = 12'h600;
			{9'd108, 8'd228}: color_data = 12'ha00;
			{9'd108, 8'd229}: color_data = 12'h900;
			{9'd108, 8'd230}: color_data = 12'h300;
			{9'd108, 8'd231}: color_data = 12'h820;
			{9'd108, 8'd232}: color_data = 12'hf30;
			{9'd108, 8'd233}: color_data = 12'hc00;
			{9'd108, 8'd234}: color_data = 12'h500;
			{9'd108, 8'd235}: color_data = 12'h200;
			{9'd108, 8'd236}: color_data = 12'h900;
			{9'd108, 8'd237}: color_data = 12'ha00;
			{9'd108, 8'd238}: color_data = 12'h700;
			{9'd108, 8'd239}: color_data = 12'h100;
			{9'd109, 8'd68}: color_data = 12'h013;
			{9'd109, 8'd69}: color_data = 12'h027;
			{9'd109, 8'd70}: color_data = 12'h016;
			{9'd109, 8'd71}: color_data = 12'h027;
			{9'd109, 8'd72}: color_data = 12'h027;
			{9'd109, 8'd73}: color_data = 12'h027;
			{9'd109, 8'd74}: color_data = 12'h027;
			{9'd109, 8'd75}: color_data = 12'h028;
			{9'd109, 8'd76}: color_data = 12'h027;
			{9'd109, 8'd77}: color_data = 12'h001;
			{9'd109, 8'd119}: color_data = 12'h000;
			{9'd109, 8'd120}: color_data = 12'h016;
			{9'd109, 8'd121}: color_data = 12'h017;
			{9'd109, 8'd122}: color_data = 12'h016;
			{9'd109, 8'd123}: color_data = 12'h027;
			{9'd109, 8'd124}: color_data = 12'h027;
			{9'd109, 8'd125}: color_data = 12'h027;
			{9'd109, 8'd126}: color_data = 12'h027;
			{9'd109, 8'd127}: color_data = 12'h028;
			{9'd109, 8'd128}: color_data = 12'h014;
			{9'd109, 8'd129}: color_data = 12'h000;
			{9'd109, 8'd170}: color_data = 12'h000;
			{9'd109, 8'd171}: color_data = 12'h002;
			{9'd109, 8'd172}: color_data = 12'h004;
			{9'd109, 8'd173}: color_data = 12'h004;
			{9'd109, 8'd174}: color_data = 12'h004;
			{9'd109, 8'd175}: color_data = 12'h004;
			{9'd109, 8'd176}: color_data = 12'h004;
			{9'd109, 8'd177}: color_data = 12'h004;
			{9'd109, 8'd178}: color_data = 12'h004;
			{9'd109, 8'd179}: color_data = 12'h004;
			{9'd109, 8'd180}: color_data = 12'h000;
			{9'd109, 8'd222}: color_data = 12'h300;
			{9'd109, 8'd223}: color_data = 12'hc30;
			{9'd109, 8'd224}: color_data = 12'hc30;
			{9'd109, 8'd225}: color_data = 12'h700;
			{9'd109, 8'd226}: color_data = 12'h100;
			{9'd109, 8'd227}: color_data = 12'h600;
			{9'd109, 8'd228}: color_data = 12'ha00;
			{9'd109, 8'd229}: color_data = 12'h900;
			{9'd109, 8'd230}: color_data = 12'h300;
			{9'd109, 8'd231}: color_data = 12'h620;
			{9'd109, 8'd232}: color_data = 12'hd40;
			{9'd109, 8'd233}: color_data = 12'ha20;
			{9'd109, 8'd234}: color_data = 12'h300;
			{9'd109, 8'd235}: color_data = 12'h200;
			{9'd109, 8'd236}: color_data = 12'h900;
			{9'd109, 8'd237}: color_data = 12'ha00;
			{9'd109, 8'd238}: color_data = 12'h700;
			{9'd109, 8'd239}: color_data = 12'h100;
			{9'd110, 8'd68}: color_data = 12'h035;
			{9'd110, 8'd69}: color_data = 12'h09e;
			{9'd110, 8'd70}: color_data = 12'h09e;
			{9'd110, 8'd71}: color_data = 12'h09e;
			{9'd110, 8'd72}: color_data = 12'h09e;
			{9'd110, 8'd73}: color_data = 12'h09e;
			{9'd110, 8'd74}: color_data = 12'h09e;
			{9'd110, 8'd75}: color_data = 12'h09e;
			{9'd110, 8'd76}: color_data = 12'h08c;
			{9'd110, 8'd77}: color_data = 12'h023;
			{9'd110, 8'd119}: color_data = 12'h000;
			{9'd110, 8'd120}: color_data = 12'h07b;
			{9'd110, 8'd121}: color_data = 12'h0ae;
			{9'd110, 8'd122}: color_data = 12'h09e;
			{9'd110, 8'd123}: color_data = 12'h09e;
			{9'd110, 8'd124}: color_data = 12'h09e;
			{9'd110, 8'd125}: color_data = 12'h09e;
			{9'd110, 8'd126}: color_data = 12'h09e;
			{9'd110, 8'd127}: color_data = 12'h09e;
			{9'd110, 8'd128}: color_data = 12'h057;
			{9'd110, 8'd129}: color_data = 12'h000;
			{9'd110, 8'd171}: color_data = 12'h000;
			{9'd110, 8'd172}: color_data = 12'h000;
			{9'd110, 8'd173}: color_data = 12'h001;
			{9'd110, 8'd174}: color_data = 12'h000;
			{9'd110, 8'd175}: color_data = 12'h000;
			{9'd110, 8'd176}: color_data = 12'h000;
			{9'd110, 8'd177}: color_data = 12'h000;
			{9'd110, 8'd178}: color_data = 12'h000;
			{9'd110, 8'd179}: color_data = 12'h000;
			{9'd110, 8'd180}: color_data = 12'h000;
			{9'd110, 8'd222}: color_data = 12'h000;
			{9'd110, 8'd223}: color_data = 12'h200;
			{9'd110, 8'd224}: color_data = 12'h300;
			{9'd110, 8'd225}: color_data = 12'h100;
			{9'd110, 8'd226}: color_data = 12'h000;
			{9'd110, 8'd227}: color_data = 12'h700;
			{9'd110, 8'd228}: color_data = 12'ha00;
			{9'd110, 8'd229}: color_data = 12'h900;
			{9'd110, 8'd230}: color_data = 12'h300;
			{9'd110, 8'd231}: color_data = 12'h100;
			{9'd110, 8'd232}: color_data = 12'h310;
			{9'd110, 8'd233}: color_data = 12'h200;
			{9'd110, 8'd234}: color_data = 12'h000;
			{9'd110, 8'd235}: color_data = 12'h300;
			{9'd110, 8'd236}: color_data = 12'h900;
			{9'd110, 8'd237}: color_data = 12'ha00;
			{9'd110, 8'd238}: color_data = 12'h700;
			{9'd110, 8'd239}: color_data = 12'h100;
			{9'd111, 8'd68}: color_data = 12'h057;
			{9'd111, 8'd69}: color_data = 12'h4ef;
			{9'd111, 8'd70}: color_data = 12'h7ef;
			{9'd111, 8'd71}: color_data = 12'h0cf;
			{9'd111, 8'd72}: color_data = 12'h0cf;
			{9'd111, 8'd73}: color_data = 12'h0df;
			{9'd111, 8'd74}: color_data = 12'h0bd;
			{9'd111, 8'd75}: color_data = 12'h068;
			{9'd111, 8'd76}: color_data = 12'h09c;
			{9'd111, 8'd77}: color_data = 12'h034;
			{9'd111, 8'd119}: color_data = 12'h000;
			{9'd111, 8'd120}: color_data = 12'h1ad;
			{9'd111, 8'd121}: color_data = 12'h8ff;
			{9'd111, 8'd122}: color_data = 12'h3df;
			{9'd111, 8'd123}: color_data = 12'h0cf;
			{9'd111, 8'd124}: color_data = 12'h0cf;
			{9'd111, 8'd125}: color_data = 12'h0cf;
			{9'd111, 8'd126}: color_data = 12'h079;
			{9'd111, 8'd127}: color_data = 12'h08b;
			{9'd111, 8'd128}: color_data = 12'h079;
			{9'd111, 8'd129}: color_data = 12'h000;
			{9'd111, 8'd222}: color_data = 12'h100;
			{9'd111, 8'd223}: color_data = 12'h400;
			{9'd111, 8'd224}: color_data = 12'h500;
			{9'd111, 8'd225}: color_data = 12'h400;
			{9'd111, 8'd226}: color_data = 12'h200;
			{9'd111, 8'd227}: color_data = 12'ha20;
			{9'd111, 8'd228}: color_data = 12'hb10;
			{9'd111, 8'd229}: color_data = 12'h900;
			{9'd111, 8'd230}: color_data = 12'h300;
			{9'd111, 8'd231}: color_data = 12'h200;
			{9'd111, 8'd232}: color_data = 12'h500;
			{9'd111, 8'd233}: color_data = 12'h500;
			{9'd111, 8'd234}: color_data = 12'h200;
			{9'd111, 8'd235}: color_data = 12'h410;
			{9'd111, 8'd236}: color_data = 12'hc20;
			{9'd111, 8'd237}: color_data = 12'ha00;
			{9'd111, 8'd238}: color_data = 12'h700;
			{9'd111, 8'd239}: color_data = 12'h100;
			{9'd112, 8'd68}: color_data = 12'h047;
			{9'd112, 8'd69}: color_data = 12'h6df;
			{9'd112, 8'd70}: color_data = 12'heff;
			{9'd112, 8'd71}: color_data = 12'h6df;
			{9'd112, 8'd72}: color_data = 12'h0bf;
			{9'd112, 8'd73}: color_data = 12'h0bf;
			{9'd112, 8'd74}: color_data = 12'h056;
			{9'd112, 8'd75}: color_data = 12'h012;
			{9'd112, 8'd76}: color_data = 12'h08b;
			{9'd112, 8'd77}: color_data = 12'h034;
			{9'd112, 8'd119}: color_data = 12'h000;
			{9'd112, 8'd120}: color_data = 12'h2ac;
			{9'd112, 8'd121}: color_data = 12'hdff;
			{9'd112, 8'd122}: color_data = 12'haef;
			{9'd112, 8'd123}: color_data = 12'h1bf;
			{9'd112, 8'd124}: color_data = 12'h0cf;
			{9'd112, 8'd125}: color_data = 12'h08b;
			{9'd112, 8'd126}: color_data = 12'h012;
			{9'd112, 8'd127}: color_data = 12'h068;
			{9'd112, 8'd128}: color_data = 12'h079;
			{9'd112, 8'd129}: color_data = 12'h000;
			{9'd112, 8'd222}: color_data = 12'h200;
			{9'd112, 8'd223}: color_data = 12'h900;
			{9'd112, 8'd224}: color_data = 12'hb00;
			{9'd112, 8'd225}: color_data = 12'h800;
			{9'd112, 8'd226}: color_data = 12'h200;
			{9'd112, 8'd227}: color_data = 12'hb30;
			{9'd112, 8'd228}: color_data = 12'hc10;
			{9'd112, 8'd229}: color_data = 12'h800;
			{9'd112, 8'd230}: color_data = 12'h300;
			{9'd112, 8'd231}: color_data = 12'h400;
			{9'd112, 8'd232}: color_data = 12'ha00;
			{9'd112, 8'd233}: color_data = 12'ha00;
			{9'd112, 8'd234}: color_data = 12'h500;
			{9'd112, 8'd235}: color_data = 12'h510;
			{9'd112, 8'd236}: color_data = 12'hd30;
			{9'd112, 8'd237}: color_data = 12'ha00;
			{9'd112, 8'd238}: color_data = 12'h700;
			{9'd112, 8'd239}: color_data = 12'h100;
			{9'd113, 8'd68}: color_data = 12'h047;
			{9'd113, 8'd69}: color_data = 12'h6df;
			{9'd113, 8'd70}: color_data = 12'hfff;
			{9'd113, 8'd71}: color_data = 12'hdff;
			{9'd113, 8'd72}: color_data = 12'h5df;
			{9'd113, 8'd73}: color_data = 12'h068;
			{9'd113, 8'd74}: color_data = 12'h000;
			{9'd113, 8'd75}: color_data = 12'h012;
			{9'd113, 8'd76}: color_data = 12'h08c;
			{9'd113, 8'd77}: color_data = 12'h034;
			{9'd113, 8'd119}: color_data = 12'h000;
			{9'd113, 8'd120}: color_data = 12'h1ac;
			{9'd113, 8'd121}: color_data = 12'hdff;
			{9'd113, 8'd122}: color_data = 12'hfff;
			{9'd113, 8'd123}: color_data = 12'h8ef;
			{9'd113, 8'd124}: color_data = 12'h19c;
			{9'd113, 8'd125}: color_data = 12'h023;
			{9'd113, 8'd127}: color_data = 12'h068;
			{9'd113, 8'd128}: color_data = 12'h079;
			{9'd113, 8'd129}: color_data = 12'h000;
			{9'd113, 8'd222}: color_data = 12'h200;
			{9'd113, 8'd223}: color_data = 12'h900;
			{9'd113, 8'd224}: color_data = 12'ha00;
			{9'd113, 8'd225}: color_data = 12'h700;
			{9'd113, 8'd226}: color_data = 12'h200;
			{9'd113, 8'd227}: color_data = 12'hb30;
			{9'd113, 8'd228}: color_data = 12'he20;
			{9'd113, 8'd229}: color_data = 12'ha00;
			{9'd113, 8'd230}: color_data = 12'h300;
			{9'd113, 8'd231}: color_data = 12'h400;
			{9'd113, 8'd232}: color_data = 12'ha00;
			{9'd113, 8'd233}: color_data = 12'ha00;
			{9'd113, 8'd234}: color_data = 12'h400;
			{9'd113, 8'd235}: color_data = 12'h510;
			{9'd113, 8'd236}: color_data = 12'hf40;
			{9'd113, 8'd237}: color_data = 12'hd10;
			{9'd113, 8'd238}: color_data = 12'h800;
			{9'd113, 8'd239}: color_data = 12'h100;
			{9'd114, 8'd68}: color_data = 12'h047;
			{9'd114, 8'd69}: color_data = 12'h6df;
			{9'd114, 8'd70}: color_data = 12'hfff;
			{9'd114, 8'd71}: color_data = 12'hfff;
			{9'd114, 8'd72}: color_data = 12'h9aa;
			{9'd114, 8'd73}: color_data = 12'h011;
			{9'd114, 8'd75}: color_data = 12'h012;
			{9'd114, 8'd76}: color_data = 12'h08c;
			{9'd114, 8'd77}: color_data = 12'h034;
			{9'd114, 8'd119}: color_data = 12'h000;
			{9'd114, 8'd120}: color_data = 12'h1ac;
			{9'd114, 8'd121}: color_data = 12'hcff;
			{9'd114, 8'd122}: color_data = 12'hfff;
			{9'd114, 8'd123}: color_data = 12'hddd;
			{9'd114, 8'd124}: color_data = 12'h345;
			{9'd114, 8'd126}: color_data = 12'h000;
			{9'd114, 8'd127}: color_data = 12'h068;
			{9'd114, 8'd128}: color_data = 12'h079;
			{9'd114, 8'd129}: color_data = 12'h000;
			{9'd114, 8'd222}: color_data = 12'h200;
			{9'd114, 8'd223}: color_data = 12'h800;
			{9'd114, 8'd224}: color_data = 12'ha00;
			{9'd114, 8'd225}: color_data = 12'h800;
			{9'd114, 8'd226}: color_data = 12'h200;
			{9'd114, 8'd227}: color_data = 12'h930;
			{9'd114, 8'd228}: color_data = 12'hd30;
			{9'd114, 8'd229}: color_data = 12'h910;
			{9'd114, 8'd230}: color_data = 12'h200;
			{9'd114, 8'd231}: color_data = 12'h400;
			{9'd114, 8'd232}: color_data = 12'h900;
			{9'd114, 8'd233}: color_data = 12'ha00;
			{9'd114, 8'd234}: color_data = 12'h400;
			{9'd114, 8'd235}: color_data = 12'h310;
			{9'd114, 8'd236}: color_data = 12'hc30;
			{9'd114, 8'd237}: color_data = 12'hc20;
			{9'd114, 8'd238}: color_data = 12'h600;
			{9'd114, 8'd239}: color_data = 12'h000;
			{9'd115, 8'd68}: color_data = 12'h047;
			{9'd115, 8'd69}: color_data = 12'h6df;
			{9'd115, 8'd70}: color_data = 12'hfff;
			{9'd115, 8'd71}: color_data = 12'hcbb;
			{9'd115, 8'd72}: color_data = 12'h323;
			{9'd115, 8'd73}: color_data = 12'h002;
			{9'd115, 8'd74}: color_data = 12'h000;
			{9'd115, 8'd75}: color_data = 12'h012;
			{9'd115, 8'd76}: color_data = 12'h08c;
			{9'd115, 8'd77}: color_data = 12'h034;
			{9'd115, 8'd119}: color_data = 12'h000;
			{9'd115, 8'd120}: color_data = 12'h1ac;
			{9'd115, 8'd121}: color_data = 12'hdff;
			{9'd115, 8'd122}: color_data = 12'hfee;
			{9'd115, 8'd123}: color_data = 12'h666;
			{9'd115, 8'd124}: color_data = 12'h002;
			{9'd115, 8'd125}: color_data = 12'h001;
			{9'd115, 8'd126}: color_data = 12'h000;
			{9'd115, 8'd127}: color_data = 12'h068;
			{9'd115, 8'd128}: color_data = 12'h079;
			{9'd115, 8'd129}: color_data = 12'h000;
			{9'd115, 8'd222}: color_data = 12'h200;
			{9'd115, 8'd223}: color_data = 12'h900;
			{9'd115, 8'd224}: color_data = 12'ha00;
			{9'd115, 8'd225}: color_data = 12'h800;
			{9'd115, 8'd226}: color_data = 12'h100;
			{9'd115, 8'd227}: color_data = 12'h100;
			{9'd115, 8'd228}: color_data = 12'h310;
			{9'd115, 8'd229}: color_data = 12'h200;
			{9'd115, 8'd230}: color_data = 12'h000;
			{9'd115, 8'd231}: color_data = 12'h500;
			{9'd115, 8'd232}: color_data = 12'ha00;
			{9'd115, 8'd233}: color_data = 12'ha00;
			{9'd115, 8'd234}: color_data = 12'h500;
			{9'd115, 8'd235}: color_data = 12'h000;
			{9'd115, 8'd236}: color_data = 12'h200;
			{9'd115, 8'd237}: color_data = 12'h300;
			{9'd115, 8'd238}: color_data = 12'h100;
			{9'd115, 8'd239}: color_data = 12'h000;
			{9'd116, 8'd68}: color_data = 12'h047;
			{9'd116, 8'd69}: color_data = 12'h6ef;
			{9'd116, 8'd70}: color_data = 12'hddc;
			{9'd116, 8'd71}: color_data = 12'h434;
			{9'd116, 8'd72}: color_data = 12'h003;
			{9'd116, 8'd73}: color_data = 12'h005;
			{9'd116, 8'd74}: color_data = 12'h002;
			{9'd116, 8'd75}: color_data = 12'h012;
			{9'd116, 8'd76}: color_data = 12'h08c;
			{9'd116, 8'd77}: color_data = 12'h034;
			{9'd116, 8'd119}: color_data = 12'h000;
			{9'd116, 8'd120}: color_data = 12'h2ad;
			{9'd116, 8'd121}: color_data = 12'hcff;
			{9'd116, 8'd122}: color_data = 12'h877;
			{9'd116, 8'd123}: color_data = 12'h002;
			{9'd116, 8'd124}: color_data = 12'h004;
			{9'd116, 8'd125}: color_data = 12'h004;
			{9'd116, 8'd126}: color_data = 12'h000;
			{9'd116, 8'd127}: color_data = 12'h068;
			{9'd116, 8'd128}: color_data = 12'h079;
			{9'd116, 8'd129}: color_data = 12'h000;
			{9'd116, 8'd222}: color_data = 12'h300;
			{9'd116, 8'd223}: color_data = 12'hc20;
			{9'd116, 8'd224}: color_data = 12'ha00;
			{9'd116, 8'd225}: color_data = 12'h800;
			{9'd116, 8'd226}: color_data = 12'h100;
			{9'd116, 8'd227}: color_data = 12'h300;
			{9'd116, 8'd228}: color_data = 12'h500;
			{9'd116, 8'd229}: color_data = 12'h500;
			{9'd116, 8'd230}: color_data = 12'h100;
			{9'd116, 8'd231}: color_data = 12'h710;
			{9'd116, 8'd232}: color_data = 12'hc10;
			{9'd116, 8'd233}: color_data = 12'h900;
			{9'd116, 8'd234}: color_data = 12'h500;
			{9'd116, 8'd235}: color_data = 12'h100;
			{9'd116, 8'd236}: color_data = 12'h500;
			{9'd116, 8'd237}: color_data = 12'h600;
			{9'd116, 8'd238}: color_data = 12'h400;
			{9'd116, 8'd239}: color_data = 12'h000;
			{9'd117, 8'd68}: color_data = 12'h057;
			{9'd117, 8'd69}: color_data = 12'h3bd;
			{9'd117, 8'd70}: color_data = 12'h555;
			{9'd117, 8'd71}: color_data = 12'h002;
			{9'd117, 8'd72}: color_data = 12'h005;
			{9'd117, 8'd73}: color_data = 12'h005;
			{9'd117, 8'd74}: color_data = 12'h004;
			{9'd117, 8'd75}: color_data = 12'h025;
			{9'd117, 8'd76}: color_data = 12'h09c;
			{9'd117, 8'd77}: color_data = 12'h034;
			{9'd117, 8'd119}: color_data = 12'h000;
			{9'd117, 8'd120}: color_data = 12'h1ac;
			{9'd117, 8'd121}: color_data = 12'h689;
			{9'd117, 8'd122}: color_data = 12'h212;
			{9'd117, 8'd123}: color_data = 12'h004;
			{9'd117, 8'd124}: color_data = 12'h005;
			{9'd117, 8'd125}: color_data = 12'h005;
			{9'd117, 8'd126}: color_data = 12'h003;
			{9'd117, 8'd127}: color_data = 12'h06a;
			{9'd117, 8'd128}: color_data = 12'h079;
			{9'd117, 8'd129}: color_data = 12'h000;
			{9'd117, 8'd222}: color_data = 12'h410;
			{9'd117, 8'd223}: color_data = 12'hd30;
			{9'd117, 8'd224}: color_data = 12'hb00;
			{9'd117, 8'd225}: color_data = 12'h700;
			{9'd117, 8'd226}: color_data = 12'h200;
			{9'd117, 8'd227}: color_data = 12'h700;
			{9'd117, 8'd228}: color_data = 12'hb00;
			{9'd117, 8'd229}: color_data = 12'ha00;
			{9'd117, 8'd230}: color_data = 12'h300;
			{9'd117, 8'd231}: color_data = 12'h820;
			{9'd117, 8'd232}: color_data = 12'hd20;
			{9'd117, 8'd233}: color_data = 12'h900;
			{9'd117, 8'd234}: color_data = 12'h500;
			{9'd117, 8'd235}: color_data = 12'h300;
			{9'd117, 8'd236}: color_data = 12'h900;
			{9'd117, 8'd237}: color_data = 12'hb00;
			{9'd117, 8'd238}: color_data = 12'h800;
			{9'd117, 8'd239}: color_data = 12'h100;
			{9'd118, 8'd68}: color_data = 12'h036;
			{9'd118, 8'd69}: color_data = 12'h047;
			{9'd118, 8'd70}: color_data = 12'h001;
			{9'd118, 8'd71}: color_data = 12'h004;
			{9'd118, 8'd72}: color_data = 12'h004;
			{9'd118, 8'd73}: color_data = 12'h004;
			{9'd118, 8'd74}: color_data = 12'h004;
			{9'd118, 8'd75}: color_data = 12'h015;
			{9'd118, 8'd76}: color_data = 12'h059;
			{9'd118, 8'd77}: color_data = 12'h023;
			{9'd118, 8'd119}: color_data = 12'h000;
			{9'd118, 8'd120}: color_data = 12'h058;
			{9'd118, 8'd121}: color_data = 12'h013;
			{9'd118, 8'd122}: color_data = 12'h002;
			{9'd118, 8'd123}: color_data = 12'h004;
			{9'd118, 8'd124}: color_data = 12'h004;
			{9'd118, 8'd125}: color_data = 12'h004;
			{9'd118, 8'd126}: color_data = 12'h004;
			{9'd118, 8'd127}: color_data = 12'h039;
			{9'd118, 8'd128}: color_data = 12'h046;
			{9'd118, 8'd129}: color_data = 12'h000;
			{9'd118, 8'd222}: color_data = 12'h410;
			{9'd118, 8'd223}: color_data = 12'he40;
			{9'd118, 8'd224}: color_data = 12'hd20;
			{9'd118, 8'd225}: color_data = 12'h800;
			{9'd118, 8'd226}: color_data = 12'h200;
			{9'd118, 8'd227}: color_data = 12'h600;
			{9'd118, 8'd228}: color_data = 12'ha00;
			{9'd118, 8'd229}: color_data = 12'h900;
			{9'd118, 8'd230}: color_data = 12'h300;
			{9'd118, 8'd231}: color_data = 12'h820;
			{9'd118, 8'd232}: color_data = 12'hf30;
			{9'd118, 8'd233}: color_data = 12'hc00;
			{9'd118, 8'd234}: color_data = 12'h500;
			{9'd118, 8'd235}: color_data = 12'h200;
			{9'd118, 8'd236}: color_data = 12'h900;
			{9'd118, 8'd237}: color_data = 12'ha00;
			{9'd118, 8'd238}: color_data = 12'h700;
			{9'd118, 8'd239}: color_data = 12'h100;
			{9'd119, 8'd68}: color_data = 12'h013;
			{9'd119, 8'd69}: color_data = 12'h027;
			{9'd119, 8'd70}: color_data = 12'h016;
			{9'd119, 8'd71}: color_data = 12'h027;
			{9'd119, 8'd72}: color_data = 12'h027;
			{9'd119, 8'd73}: color_data = 12'h027;
			{9'd119, 8'd74}: color_data = 12'h027;
			{9'd119, 8'd75}: color_data = 12'h028;
			{9'd119, 8'd76}: color_data = 12'h027;
			{9'd119, 8'd77}: color_data = 12'h001;
			{9'd119, 8'd119}: color_data = 12'h000;
			{9'd119, 8'd120}: color_data = 12'h016;
			{9'd119, 8'd121}: color_data = 12'h017;
			{9'd119, 8'd122}: color_data = 12'h016;
			{9'd119, 8'd123}: color_data = 12'h027;
			{9'd119, 8'd124}: color_data = 12'h027;
			{9'd119, 8'd125}: color_data = 12'h027;
			{9'd119, 8'd126}: color_data = 12'h027;
			{9'd119, 8'd127}: color_data = 12'h028;
			{9'd119, 8'd128}: color_data = 12'h014;
			{9'd119, 8'd129}: color_data = 12'h000;
			{9'd119, 8'd222}: color_data = 12'h300;
			{9'd119, 8'd223}: color_data = 12'hc30;
			{9'd119, 8'd224}: color_data = 12'hc30;
			{9'd119, 8'd225}: color_data = 12'h700;
			{9'd119, 8'd226}: color_data = 12'h100;
			{9'd119, 8'd227}: color_data = 12'h600;
			{9'd119, 8'd228}: color_data = 12'ha00;
			{9'd119, 8'd229}: color_data = 12'h900;
			{9'd119, 8'd230}: color_data = 12'h300;
			{9'd119, 8'd231}: color_data = 12'h620;
			{9'd119, 8'd232}: color_data = 12'hd40;
			{9'd119, 8'd233}: color_data = 12'ha20;
			{9'd119, 8'd234}: color_data = 12'h300;
			{9'd119, 8'd235}: color_data = 12'h200;
			{9'd119, 8'd236}: color_data = 12'h800;
			{9'd119, 8'd237}: color_data = 12'ha00;
			{9'd119, 8'd238}: color_data = 12'h700;
			{9'd119, 8'd239}: color_data = 12'h100;
			{9'd120, 8'd68}: color_data = 12'h035;
			{9'd120, 8'd69}: color_data = 12'h09e;
			{9'd120, 8'd70}: color_data = 12'h09e;
			{9'd120, 8'd71}: color_data = 12'h09e;
			{9'd120, 8'd72}: color_data = 12'h09e;
			{9'd120, 8'd73}: color_data = 12'h09e;
			{9'd120, 8'd74}: color_data = 12'h09e;
			{9'd120, 8'd75}: color_data = 12'h09e;
			{9'd120, 8'd76}: color_data = 12'h08c;
			{9'd120, 8'd77}: color_data = 12'h023;
			{9'd120, 8'd119}: color_data = 12'h000;
			{9'd120, 8'd120}: color_data = 12'h07b;
			{9'd120, 8'd121}: color_data = 12'h0ae;
			{9'd120, 8'd122}: color_data = 12'h09e;
			{9'd120, 8'd123}: color_data = 12'h09e;
			{9'd120, 8'd124}: color_data = 12'h09e;
			{9'd120, 8'd125}: color_data = 12'h09e;
			{9'd120, 8'd126}: color_data = 12'h09e;
			{9'd120, 8'd127}: color_data = 12'h09e;
			{9'd120, 8'd128}: color_data = 12'h057;
			{9'd120, 8'd129}: color_data = 12'h000;
			{9'd120, 8'd222}: color_data = 12'h000;
			{9'd120, 8'd223}: color_data = 12'h200;
			{9'd120, 8'd224}: color_data = 12'h300;
			{9'd120, 8'd225}: color_data = 12'h100;
			{9'd120, 8'd226}: color_data = 12'h000;
			{9'd120, 8'd227}: color_data = 12'h700;
			{9'd120, 8'd228}: color_data = 12'ha00;
			{9'd120, 8'd229}: color_data = 12'h900;
			{9'd120, 8'd230}: color_data = 12'h300;
			{9'd120, 8'd231}: color_data = 12'h100;
			{9'd120, 8'd232}: color_data = 12'h310;
			{9'd120, 8'd233}: color_data = 12'h200;
			{9'd120, 8'd234}: color_data = 12'h000;
			{9'd120, 8'd235}: color_data = 12'h300;
			{9'd120, 8'd236}: color_data = 12'h900;
			{9'd120, 8'd237}: color_data = 12'ha00;
			{9'd120, 8'd238}: color_data = 12'h700;
			{9'd120, 8'd239}: color_data = 12'h100;
			{9'd121, 8'd68}: color_data = 12'h057;
			{9'd121, 8'd69}: color_data = 12'h4ef;
			{9'd121, 8'd70}: color_data = 12'h7ef;
			{9'd121, 8'd71}: color_data = 12'h0cf;
			{9'd121, 8'd72}: color_data = 12'h0cf;
			{9'd121, 8'd73}: color_data = 12'h0df;
			{9'd121, 8'd74}: color_data = 12'h0bd;
			{9'd121, 8'd75}: color_data = 12'h068;
			{9'd121, 8'd76}: color_data = 12'h09c;
			{9'd121, 8'd77}: color_data = 12'h034;
			{9'd121, 8'd119}: color_data = 12'h000;
			{9'd121, 8'd120}: color_data = 12'h1ad;
			{9'd121, 8'd121}: color_data = 12'h8ff;
			{9'd121, 8'd122}: color_data = 12'h3df;
			{9'd121, 8'd123}: color_data = 12'h0cf;
			{9'd121, 8'd124}: color_data = 12'h0cf;
			{9'd121, 8'd125}: color_data = 12'h0cf;
			{9'd121, 8'd126}: color_data = 12'h07a;
			{9'd121, 8'd127}: color_data = 12'h08b;
			{9'd121, 8'd128}: color_data = 12'h079;
			{9'd121, 8'd129}: color_data = 12'h000;
			{9'd121, 8'd222}: color_data = 12'h100;
			{9'd121, 8'd223}: color_data = 12'h400;
			{9'd121, 8'd224}: color_data = 12'h500;
			{9'd121, 8'd225}: color_data = 12'h400;
			{9'd121, 8'd226}: color_data = 12'h200;
			{9'd121, 8'd227}: color_data = 12'ha20;
			{9'd121, 8'd228}: color_data = 12'hb10;
			{9'd121, 8'd229}: color_data = 12'h900;
			{9'd121, 8'd230}: color_data = 12'h300;
			{9'd121, 8'd231}: color_data = 12'h200;
			{9'd121, 8'd232}: color_data = 12'h500;
			{9'd121, 8'd233}: color_data = 12'h500;
			{9'd121, 8'd234}: color_data = 12'h200;
			{9'd121, 8'd235}: color_data = 12'h410;
			{9'd121, 8'd236}: color_data = 12'hc20;
			{9'd121, 8'd237}: color_data = 12'ha00;
			{9'd121, 8'd238}: color_data = 12'h700;
			{9'd121, 8'd239}: color_data = 12'h100;
			{9'd122, 8'd68}: color_data = 12'h047;
			{9'd122, 8'd69}: color_data = 12'h6df;
			{9'd122, 8'd70}: color_data = 12'heff;
			{9'd122, 8'd71}: color_data = 12'h6df;
			{9'd122, 8'd72}: color_data = 12'h0bf;
			{9'd122, 8'd73}: color_data = 12'h0be;
			{9'd122, 8'd74}: color_data = 12'h056;
			{9'd122, 8'd75}: color_data = 12'h012;
			{9'd122, 8'd76}: color_data = 12'h08b;
			{9'd122, 8'd77}: color_data = 12'h034;
			{9'd122, 8'd119}: color_data = 12'h000;
			{9'd122, 8'd120}: color_data = 12'h2ac;
			{9'd122, 8'd121}: color_data = 12'hdff;
			{9'd122, 8'd122}: color_data = 12'haef;
			{9'd122, 8'd123}: color_data = 12'h1bf;
			{9'd122, 8'd124}: color_data = 12'h0cf;
			{9'd122, 8'd125}: color_data = 12'h08b;
			{9'd122, 8'd126}: color_data = 12'h012;
			{9'd122, 8'd127}: color_data = 12'h068;
			{9'd122, 8'd128}: color_data = 12'h079;
			{9'd122, 8'd129}: color_data = 12'h000;
			{9'd122, 8'd222}: color_data = 12'h200;
			{9'd122, 8'd223}: color_data = 12'h900;
			{9'd122, 8'd224}: color_data = 12'hb00;
			{9'd122, 8'd225}: color_data = 12'h800;
			{9'd122, 8'd226}: color_data = 12'h200;
			{9'd122, 8'd227}: color_data = 12'hb30;
			{9'd122, 8'd228}: color_data = 12'hc10;
			{9'd122, 8'd229}: color_data = 12'h800;
			{9'd122, 8'd230}: color_data = 12'h300;
			{9'd122, 8'd231}: color_data = 12'h400;
			{9'd122, 8'd232}: color_data = 12'ha00;
			{9'd122, 8'd233}: color_data = 12'ha00;
			{9'd122, 8'd234}: color_data = 12'h500;
			{9'd122, 8'd235}: color_data = 12'h510;
			{9'd122, 8'd236}: color_data = 12'hd30;
			{9'd122, 8'd237}: color_data = 12'ha00;
			{9'd122, 8'd238}: color_data = 12'h700;
			{9'd122, 8'd239}: color_data = 12'h100;
			{9'd123, 8'd68}: color_data = 12'h047;
			{9'd123, 8'd69}: color_data = 12'h6df;
			{9'd123, 8'd70}: color_data = 12'hfff;
			{9'd123, 8'd71}: color_data = 12'hdff;
			{9'd123, 8'd72}: color_data = 12'h5df;
			{9'd123, 8'd73}: color_data = 12'h068;
			{9'd123, 8'd74}: color_data = 12'h000;
			{9'd123, 8'd75}: color_data = 12'h012;
			{9'd123, 8'd76}: color_data = 12'h08c;
			{9'd123, 8'd77}: color_data = 12'h034;
			{9'd123, 8'd119}: color_data = 12'h000;
			{9'd123, 8'd120}: color_data = 12'h1ac;
			{9'd123, 8'd121}: color_data = 12'hdff;
			{9'd123, 8'd122}: color_data = 12'hfff;
			{9'd123, 8'd123}: color_data = 12'h8ef;
			{9'd123, 8'd124}: color_data = 12'h19c;
			{9'd123, 8'd125}: color_data = 12'h023;
			{9'd123, 8'd127}: color_data = 12'h068;
			{9'd123, 8'd128}: color_data = 12'h079;
			{9'd123, 8'd129}: color_data = 12'h000;
			{9'd123, 8'd222}: color_data = 12'h200;
			{9'd123, 8'd223}: color_data = 12'h900;
			{9'd123, 8'd224}: color_data = 12'ha00;
			{9'd123, 8'd225}: color_data = 12'h700;
			{9'd123, 8'd226}: color_data = 12'h200;
			{9'd123, 8'd227}: color_data = 12'hb30;
			{9'd123, 8'd228}: color_data = 12'he20;
			{9'd123, 8'd229}: color_data = 12'ha00;
			{9'd123, 8'd230}: color_data = 12'h300;
			{9'd123, 8'd231}: color_data = 12'h400;
			{9'd123, 8'd232}: color_data = 12'ha00;
			{9'd123, 8'd233}: color_data = 12'ha00;
			{9'd123, 8'd234}: color_data = 12'h400;
			{9'd123, 8'd235}: color_data = 12'h510;
			{9'd123, 8'd236}: color_data = 12'hf40;
			{9'd123, 8'd237}: color_data = 12'hd10;
			{9'd123, 8'd238}: color_data = 12'h800;
			{9'd123, 8'd239}: color_data = 12'h100;
			{9'd124, 8'd68}: color_data = 12'h047;
			{9'd124, 8'd69}: color_data = 12'h6df;
			{9'd124, 8'd70}: color_data = 12'hfff;
			{9'd124, 8'd71}: color_data = 12'hfff;
			{9'd124, 8'd72}: color_data = 12'h9aa;
			{9'd124, 8'd73}: color_data = 12'h011;
			{9'd124, 8'd75}: color_data = 12'h012;
			{9'd124, 8'd76}: color_data = 12'h08c;
			{9'd124, 8'd77}: color_data = 12'h034;
			{9'd124, 8'd119}: color_data = 12'h000;
			{9'd124, 8'd120}: color_data = 12'h1ac;
			{9'd124, 8'd121}: color_data = 12'hcff;
			{9'd124, 8'd122}: color_data = 12'hfff;
			{9'd124, 8'd123}: color_data = 12'hddd;
			{9'd124, 8'd124}: color_data = 12'h345;
			{9'd124, 8'd126}: color_data = 12'h000;
			{9'd124, 8'd127}: color_data = 12'h068;
			{9'd124, 8'd128}: color_data = 12'h079;
			{9'd124, 8'd129}: color_data = 12'h000;
			{9'd124, 8'd222}: color_data = 12'h200;
			{9'd124, 8'd223}: color_data = 12'h800;
			{9'd124, 8'd224}: color_data = 12'ha00;
			{9'd124, 8'd225}: color_data = 12'h700;
			{9'd124, 8'd226}: color_data = 12'h200;
			{9'd124, 8'd227}: color_data = 12'h920;
			{9'd124, 8'd228}: color_data = 12'hd30;
			{9'd124, 8'd229}: color_data = 12'h910;
			{9'd124, 8'd230}: color_data = 12'h200;
			{9'd124, 8'd231}: color_data = 12'h400;
			{9'd124, 8'd232}: color_data = 12'h900;
			{9'd124, 8'd233}: color_data = 12'ha00;
			{9'd124, 8'd234}: color_data = 12'h400;
			{9'd124, 8'd235}: color_data = 12'h310;
			{9'd124, 8'd236}: color_data = 12'hc30;
			{9'd124, 8'd237}: color_data = 12'hc20;
			{9'd124, 8'd238}: color_data = 12'h600;
			{9'd124, 8'd239}: color_data = 12'h000;
			{9'd125, 8'd68}: color_data = 12'h047;
			{9'd125, 8'd69}: color_data = 12'h6df;
			{9'd125, 8'd70}: color_data = 12'hfff;
			{9'd125, 8'd71}: color_data = 12'hcbb;
			{9'd125, 8'd72}: color_data = 12'h323;
			{9'd125, 8'd73}: color_data = 12'h002;
			{9'd125, 8'd74}: color_data = 12'h000;
			{9'd125, 8'd75}: color_data = 12'h012;
			{9'd125, 8'd76}: color_data = 12'h08c;
			{9'd125, 8'd77}: color_data = 12'h034;
			{9'd125, 8'd119}: color_data = 12'h000;
			{9'd125, 8'd120}: color_data = 12'h1ac;
			{9'd125, 8'd121}: color_data = 12'hdff;
			{9'd125, 8'd122}: color_data = 12'hfee;
			{9'd125, 8'd123}: color_data = 12'h666;
			{9'd125, 8'd124}: color_data = 12'h002;
			{9'd125, 8'd125}: color_data = 12'h001;
			{9'd125, 8'd126}: color_data = 12'h000;
			{9'd125, 8'd127}: color_data = 12'h068;
			{9'd125, 8'd128}: color_data = 12'h079;
			{9'd125, 8'd129}: color_data = 12'h000;
			{9'd125, 8'd222}: color_data = 12'h200;
			{9'd125, 8'd223}: color_data = 12'h900;
			{9'd125, 8'd224}: color_data = 12'ha00;
			{9'd125, 8'd225}: color_data = 12'h800;
			{9'd125, 8'd226}: color_data = 12'h100;
			{9'd125, 8'd227}: color_data = 12'h100;
			{9'd125, 8'd228}: color_data = 12'h310;
			{9'd125, 8'd229}: color_data = 12'h200;
			{9'd125, 8'd230}: color_data = 12'h000;
			{9'd125, 8'd231}: color_data = 12'h500;
			{9'd125, 8'd232}: color_data = 12'ha00;
			{9'd125, 8'd233}: color_data = 12'ha00;
			{9'd125, 8'd234}: color_data = 12'h500;
			{9'd125, 8'd235}: color_data = 12'h000;
			{9'd125, 8'd236}: color_data = 12'h200;
			{9'd125, 8'd237}: color_data = 12'h300;
			{9'd125, 8'd238}: color_data = 12'h100;
			{9'd125, 8'd239}: color_data = 12'h000;
			{9'd126, 8'd68}: color_data = 12'h047;
			{9'd126, 8'd69}: color_data = 12'h6ef;
			{9'd126, 8'd70}: color_data = 12'hddc;
			{9'd126, 8'd71}: color_data = 12'h434;
			{9'd126, 8'd72}: color_data = 12'h003;
			{9'd126, 8'd73}: color_data = 12'h005;
			{9'd126, 8'd74}: color_data = 12'h002;
			{9'd126, 8'd75}: color_data = 12'h012;
			{9'd126, 8'd76}: color_data = 12'h08c;
			{9'd126, 8'd77}: color_data = 12'h034;
			{9'd126, 8'd119}: color_data = 12'h000;
			{9'd126, 8'd120}: color_data = 12'h2ad;
			{9'd126, 8'd121}: color_data = 12'hcff;
			{9'd126, 8'd122}: color_data = 12'h877;
			{9'd126, 8'd123}: color_data = 12'h002;
			{9'd126, 8'd124}: color_data = 12'h004;
			{9'd126, 8'd125}: color_data = 12'h004;
			{9'd126, 8'd126}: color_data = 12'h000;
			{9'd126, 8'd127}: color_data = 12'h068;
			{9'd126, 8'd128}: color_data = 12'h079;
			{9'd126, 8'd129}: color_data = 12'h000;
			{9'd126, 8'd222}: color_data = 12'h300;
			{9'd126, 8'd223}: color_data = 12'hc20;
			{9'd126, 8'd224}: color_data = 12'ha00;
			{9'd126, 8'd225}: color_data = 12'h800;
			{9'd126, 8'd226}: color_data = 12'h100;
			{9'd126, 8'd227}: color_data = 12'h300;
			{9'd126, 8'd228}: color_data = 12'h500;
			{9'd126, 8'd229}: color_data = 12'h500;
			{9'd126, 8'd230}: color_data = 12'h100;
			{9'd126, 8'd231}: color_data = 12'h710;
			{9'd126, 8'd232}: color_data = 12'hc10;
			{9'd126, 8'd233}: color_data = 12'h900;
			{9'd126, 8'd234}: color_data = 12'h500;
			{9'd126, 8'd235}: color_data = 12'h100;
			{9'd126, 8'd236}: color_data = 12'h500;
			{9'd126, 8'd237}: color_data = 12'h500;
			{9'd126, 8'd238}: color_data = 12'h400;
			{9'd126, 8'd239}: color_data = 12'h000;
			{9'd127, 8'd68}: color_data = 12'h057;
			{9'd127, 8'd69}: color_data = 12'h3bd;
			{9'd127, 8'd70}: color_data = 12'h555;
			{9'd127, 8'd71}: color_data = 12'h002;
			{9'd127, 8'd72}: color_data = 12'h005;
			{9'd127, 8'd73}: color_data = 12'h005;
			{9'd127, 8'd74}: color_data = 12'h004;
			{9'd127, 8'd75}: color_data = 12'h025;
			{9'd127, 8'd76}: color_data = 12'h09c;
			{9'd127, 8'd77}: color_data = 12'h034;
			{9'd127, 8'd119}: color_data = 12'h000;
			{9'd127, 8'd120}: color_data = 12'h1ac;
			{9'd127, 8'd121}: color_data = 12'h689;
			{9'd127, 8'd122}: color_data = 12'h212;
			{9'd127, 8'd123}: color_data = 12'h004;
			{9'd127, 8'd124}: color_data = 12'h005;
			{9'd127, 8'd125}: color_data = 12'h005;
			{9'd127, 8'd126}: color_data = 12'h003;
			{9'd127, 8'd127}: color_data = 12'h06a;
			{9'd127, 8'd128}: color_data = 12'h079;
			{9'd127, 8'd129}: color_data = 12'h000;
			{9'd127, 8'd222}: color_data = 12'h410;
			{9'd127, 8'd223}: color_data = 12'hd30;
			{9'd127, 8'd224}: color_data = 12'hb00;
			{9'd127, 8'd225}: color_data = 12'h700;
			{9'd127, 8'd226}: color_data = 12'h200;
			{9'd127, 8'd227}: color_data = 12'h700;
			{9'd127, 8'd228}: color_data = 12'hb00;
			{9'd127, 8'd229}: color_data = 12'ha00;
			{9'd127, 8'd230}: color_data = 12'h300;
			{9'd127, 8'd231}: color_data = 12'h820;
			{9'd127, 8'd232}: color_data = 12'hd20;
			{9'd127, 8'd233}: color_data = 12'h900;
			{9'd127, 8'd234}: color_data = 12'h500;
			{9'd127, 8'd235}: color_data = 12'h300;
			{9'd127, 8'd236}: color_data = 12'h900;
			{9'd127, 8'd237}: color_data = 12'hb00;
			{9'd127, 8'd238}: color_data = 12'h800;
			{9'd127, 8'd239}: color_data = 12'h100;
			{9'd128, 8'd68}: color_data = 12'h035;
			{9'd128, 8'd69}: color_data = 12'h047;
			{9'd128, 8'd70}: color_data = 12'h001;
			{9'd128, 8'd71}: color_data = 12'h004;
			{9'd128, 8'd72}: color_data = 12'h004;
			{9'd128, 8'd73}: color_data = 12'h004;
			{9'd128, 8'd74}: color_data = 12'h004;
			{9'd128, 8'd75}: color_data = 12'h015;
			{9'd128, 8'd76}: color_data = 12'h059;
			{9'd128, 8'd77}: color_data = 12'h023;
			{9'd128, 8'd119}: color_data = 12'h000;
			{9'd128, 8'd120}: color_data = 12'h058;
			{9'd128, 8'd121}: color_data = 12'h013;
			{9'd128, 8'd122}: color_data = 12'h002;
			{9'd128, 8'd123}: color_data = 12'h004;
			{9'd128, 8'd124}: color_data = 12'h004;
			{9'd128, 8'd125}: color_data = 12'h004;
			{9'd128, 8'd126}: color_data = 12'h004;
			{9'd128, 8'd127}: color_data = 12'h038;
			{9'd128, 8'd128}: color_data = 12'h046;
			{9'd128, 8'd129}: color_data = 12'h000;
			{9'd128, 8'd222}: color_data = 12'h410;
			{9'd128, 8'd223}: color_data = 12'he40;
			{9'd128, 8'd224}: color_data = 12'hd20;
			{9'd128, 8'd225}: color_data = 12'h800;
			{9'd128, 8'd226}: color_data = 12'h200;
			{9'd128, 8'd227}: color_data = 12'h600;
			{9'd128, 8'd228}: color_data = 12'ha00;
			{9'd128, 8'd229}: color_data = 12'h900;
			{9'd128, 8'd230}: color_data = 12'h300;
			{9'd128, 8'd231}: color_data = 12'h820;
			{9'd128, 8'd232}: color_data = 12'hf30;
			{9'd128, 8'd233}: color_data = 12'hc00;
			{9'd128, 8'd234}: color_data = 12'h500;
			{9'd128, 8'd235}: color_data = 12'h200;
			{9'd128, 8'd236}: color_data = 12'h900;
			{9'd128, 8'd237}: color_data = 12'ha00;
			{9'd128, 8'd238}: color_data = 12'h700;
			{9'd128, 8'd239}: color_data = 12'h100;
			{9'd129, 8'd68}: color_data = 12'h013;
			{9'd129, 8'd69}: color_data = 12'h027;
			{9'd129, 8'd70}: color_data = 12'h016;
			{9'd129, 8'd71}: color_data = 12'h027;
			{9'd129, 8'd72}: color_data = 12'h027;
			{9'd129, 8'd73}: color_data = 12'h027;
			{9'd129, 8'd74}: color_data = 12'h027;
			{9'd129, 8'd75}: color_data = 12'h028;
			{9'd129, 8'd76}: color_data = 12'h027;
			{9'd129, 8'd77}: color_data = 12'h001;
			{9'd129, 8'd119}: color_data = 12'h000;
			{9'd129, 8'd120}: color_data = 12'h016;
			{9'd129, 8'd121}: color_data = 12'h017;
			{9'd129, 8'd122}: color_data = 12'h016;
			{9'd129, 8'd123}: color_data = 12'h027;
			{9'd129, 8'd124}: color_data = 12'h027;
			{9'd129, 8'd125}: color_data = 12'h027;
			{9'd129, 8'd126}: color_data = 12'h027;
			{9'd129, 8'd127}: color_data = 12'h028;
			{9'd129, 8'd128}: color_data = 12'h014;
			{9'd129, 8'd129}: color_data = 12'h000;
			{9'd129, 8'd222}: color_data = 12'h300;
			{9'd129, 8'd223}: color_data = 12'hc30;
			{9'd129, 8'd224}: color_data = 12'hc30;
			{9'd129, 8'd225}: color_data = 12'h600;
			{9'd129, 8'd226}: color_data = 12'h100;
			{9'd129, 8'd227}: color_data = 12'h600;
			{9'd129, 8'd228}: color_data = 12'ha00;
			{9'd129, 8'd229}: color_data = 12'h900;
			{9'd129, 8'd230}: color_data = 12'h300;
			{9'd129, 8'd231}: color_data = 12'h620;
			{9'd129, 8'd232}: color_data = 12'hd40;
			{9'd129, 8'd233}: color_data = 12'ha20;
			{9'd129, 8'd234}: color_data = 12'h300;
			{9'd129, 8'd235}: color_data = 12'h200;
			{9'd129, 8'd236}: color_data = 12'h900;
			{9'd129, 8'd237}: color_data = 12'ha00;
			{9'd129, 8'd238}: color_data = 12'h700;
			{9'd129, 8'd239}: color_data = 12'h100;
			{9'd130, 8'd68}: color_data = 12'h035;
			{9'd130, 8'd69}: color_data = 12'h09e;
			{9'd130, 8'd70}: color_data = 12'h09e;
			{9'd130, 8'd71}: color_data = 12'h09e;
			{9'd130, 8'd72}: color_data = 12'h09e;
			{9'd130, 8'd73}: color_data = 12'h09e;
			{9'd130, 8'd74}: color_data = 12'h09e;
			{9'd130, 8'd75}: color_data = 12'h09e;
			{9'd130, 8'd76}: color_data = 12'h08c;
			{9'd130, 8'd77}: color_data = 12'h023;
			{9'd130, 8'd119}: color_data = 12'h000;
			{9'd130, 8'd120}: color_data = 12'h07b;
			{9'd130, 8'd121}: color_data = 12'h0ae;
			{9'd130, 8'd122}: color_data = 12'h09e;
			{9'd130, 8'd123}: color_data = 12'h09e;
			{9'd130, 8'd124}: color_data = 12'h09e;
			{9'd130, 8'd125}: color_data = 12'h09e;
			{9'd130, 8'd126}: color_data = 12'h09e;
			{9'd130, 8'd127}: color_data = 12'h09e;
			{9'd130, 8'd128}: color_data = 12'h057;
			{9'd130, 8'd129}: color_data = 12'h000;
			{9'd130, 8'd222}: color_data = 12'h000;
			{9'd130, 8'd223}: color_data = 12'h200;
			{9'd130, 8'd224}: color_data = 12'h300;
			{9'd130, 8'd225}: color_data = 12'h100;
			{9'd130, 8'd226}: color_data = 12'h000;
			{9'd130, 8'd227}: color_data = 12'h700;
			{9'd130, 8'd228}: color_data = 12'ha00;
			{9'd130, 8'd229}: color_data = 12'h900;
			{9'd130, 8'd230}: color_data = 12'h300;
			{9'd130, 8'd231}: color_data = 12'h100;
			{9'd130, 8'd232}: color_data = 12'h300;
			{9'd130, 8'd233}: color_data = 12'h200;
			{9'd130, 8'd234}: color_data = 12'h000;
			{9'd130, 8'd235}: color_data = 12'h300;
			{9'd130, 8'd236}: color_data = 12'h900;
			{9'd130, 8'd237}: color_data = 12'ha00;
			{9'd130, 8'd238}: color_data = 12'h700;
			{9'd130, 8'd239}: color_data = 12'h100;
			{9'd131, 8'd68}: color_data = 12'h057;
			{9'd131, 8'd69}: color_data = 12'h4ef;
			{9'd131, 8'd70}: color_data = 12'h7ef;
			{9'd131, 8'd71}: color_data = 12'h0cf;
			{9'd131, 8'd72}: color_data = 12'h0cf;
			{9'd131, 8'd73}: color_data = 12'h0df;
			{9'd131, 8'd74}: color_data = 12'h0bd;
			{9'd131, 8'd75}: color_data = 12'h068;
			{9'd131, 8'd76}: color_data = 12'h09c;
			{9'd131, 8'd77}: color_data = 12'h034;
			{9'd131, 8'd119}: color_data = 12'h000;
			{9'd131, 8'd120}: color_data = 12'h1ad;
			{9'd131, 8'd121}: color_data = 12'h8ff;
			{9'd131, 8'd122}: color_data = 12'h3df;
			{9'd131, 8'd123}: color_data = 12'h0cf;
			{9'd131, 8'd124}: color_data = 12'h0cf;
			{9'd131, 8'd125}: color_data = 12'h0cf;
			{9'd131, 8'd126}: color_data = 12'h079;
			{9'd131, 8'd127}: color_data = 12'h08b;
			{9'd131, 8'd128}: color_data = 12'h079;
			{9'd131, 8'd129}: color_data = 12'h000;
			{9'd131, 8'd222}: color_data = 12'h100;
			{9'd131, 8'd223}: color_data = 12'h400;
			{9'd131, 8'd224}: color_data = 12'h500;
			{9'd131, 8'd225}: color_data = 12'h400;
			{9'd131, 8'd226}: color_data = 12'h200;
			{9'd131, 8'd227}: color_data = 12'ha20;
			{9'd131, 8'd228}: color_data = 12'hb10;
			{9'd131, 8'd229}: color_data = 12'h900;
			{9'd131, 8'd230}: color_data = 12'h300;
			{9'd131, 8'd231}: color_data = 12'h200;
			{9'd131, 8'd232}: color_data = 12'h500;
			{9'd131, 8'd233}: color_data = 12'h500;
			{9'd131, 8'd234}: color_data = 12'h200;
			{9'd131, 8'd235}: color_data = 12'h410;
			{9'd131, 8'd236}: color_data = 12'hc20;
			{9'd131, 8'd237}: color_data = 12'ha00;
			{9'd131, 8'd238}: color_data = 12'h700;
			{9'd131, 8'd239}: color_data = 12'h100;
			{9'd132, 8'd68}: color_data = 12'h047;
			{9'd132, 8'd69}: color_data = 12'h6df;
			{9'd132, 8'd70}: color_data = 12'heff;
			{9'd132, 8'd71}: color_data = 12'h6df;
			{9'd132, 8'd72}: color_data = 12'h0bf;
			{9'd132, 8'd73}: color_data = 12'h0be;
			{9'd132, 8'd74}: color_data = 12'h056;
			{9'd132, 8'd75}: color_data = 12'h012;
			{9'd132, 8'd76}: color_data = 12'h08b;
			{9'd132, 8'd77}: color_data = 12'h034;
			{9'd132, 8'd119}: color_data = 12'h000;
			{9'd132, 8'd120}: color_data = 12'h2ac;
			{9'd132, 8'd121}: color_data = 12'hdff;
			{9'd132, 8'd122}: color_data = 12'haef;
			{9'd132, 8'd123}: color_data = 12'h1cf;
			{9'd132, 8'd124}: color_data = 12'h0cf;
			{9'd132, 8'd125}: color_data = 12'h08b;
			{9'd132, 8'd126}: color_data = 12'h012;
			{9'd132, 8'd127}: color_data = 12'h068;
			{9'd132, 8'd128}: color_data = 12'h079;
			{9'd132, 8'd129}: color_data = 12'h000;
			{9'd132, 8'd222}: color_data = 12'h200;
			{9'd132, 8'd223}: color_data = 12'h900;
			{9'd132, 8'd224}: color_data = 12'hb00;
			{9'd132, 8'd225}: color_data = 12'h800;
			{9'd132, 8'd226}: color_data = 12'h200;
			{9'd132, 8'd227}: color_data = 12'hb30;
			{9'd132, 8'd228}: color_data = 12'hc10;
			{9'd132, 8'd229}: color_data = 12'h800;
			{9'd132, 8'd230}: color_data = 12'h300;
			{9'd132, 8'd231}: color_data = 12'h500;
			{9'd132, 8'd232}: color_data = 12'ha00;
			{9'd132, 8'd233}: color_data = 12'ha00;
			{9'd132, 8'd234}: color_data = 12'h500;
			{9'd132, 8'd235}: color_data = 12'h510;
			{9'd132, 8'd236}: color_data = 12'hd30;
			{9'd132, 8'd237}: color_data = 12'ha00;
			{9'd132, 8'd238}: color_data = 12'h700;
			{9'd132, 8'd239}: color_data = 12'h100;
			{9'd133, 8'd68}: color_data = 12'h047;
			{9'd133, 8'd69}: color_data = 12'h6df;
			{9'd133, 8'd70}: color_data = 12'hfff;
			{9'd133, 8'd71}: color_data = 12'hdff;
			{9'd133, 8'd72}: color_data = 12'h5df;
			{9'd133, 8'd73}: color_data = 12'h068;
			{9'd133, 8'd74}: color_data = 12'h000;
			{9'd133, 8'd75}: color_data = 12'h012;
			{9'd133, 8'd76}: color_data = 12'h08c;
			{9'd133, 8'd77}: color_data = 12'h034;
			{9'd133, 8'd119}: color_data = 12'h000;
			{9'd133, 8'd120}: color_data = 12'h1ac;
			{9'd133, 8'd121}: color_data = 12'hdff;
			{9'd133, 8'd122}: color_data = 12'hfff;
			{9'd133, 8'd123}: color_data = 12'h9ef;
			{9'd133, 8'd124}: color_data = 12'h19c;
			{9'd133, 8'd125}: color_data = 12'h023;
			{9'd133, 8'd127}: color_data = 12'h068;
			{9'd133, 8'd128}: color_data = 12'h079;
			{9'd133, 8'd129}: color_data = 12'h000;
			{9'd133, 8'd222}: color_data = 12'h200;
			{9'd133, 8'd223}: color_data = 12'h900;
			{9'd133, 8'd224}: color_data = 12'ha00;
			{9'd133, 8'd225}: color_data = 12'h700;
			{9'd133, 8'd226}: color_data = 12'h200;
			{9'd133, 8'd227}: color_data = 12'hb30;
			{9'd133, 8'd228}: color_data = 12'he20;
			{9'd133, 8'd229}: color_data = 12'ha00;
			{9'd133, 8'd230}: color_data = 12'h300;
			{9'd133, 8'd231}: color_data = 12'h400;
			{9'd133, 8'd232}: color_data = 12'ha00;
			{9'd133, 8'd233}: color_data = 12'ha00;
			{9'd133, 8'd234}: color_data = 12'h400;
			{9'd133, 8'd235}: color_data = 12'h510;
			{9'd133, 8'd236}: color_data = 12'hf40;
			{9'd133, 8'd237}: color_data = 12'hd10;
			{9'd133, 8'd238}: color_data = 12'h800;
			{9'd133, 8'd239}: color_data = 12'h100;
			{9'd134, 8'd68}: color_data = 12'h047;
			{9'd134, 8'd69}: color_data = 12'h6df;
			{9'd134, 8'd70}: color_data = 12'hfff;
			{9'd134, 8'd71}: color_data = 12'hfff;
			{9'd134, 8'd72}: color_data = 12'h9aa;
			{9'd134, 8'd73}: color_data = 12'h011;
			{9'd134, 8'd75}: color_data = 12'h012;
			{9'd134, 8'd76}: color_data = 12'h08c;
			{9'd134, 8'd77}: color_data = 12'h034;
			{9'd134, 8'd119}: color_data = 12'h000;
			{9'd134, 8'd120}: color_data = 12'h1ac;
			{9'd134, 8'd121}: color_data = 12'hcff;
			{9'd134, 8'd122}: color_data = 12'hfff;
			{9'd134, 8'd123}: color_data = 12'hddd;
			{9'd134, 8'd124}: color_data = 12'h345;
			{9'd134, 8'd126}: color_data = 12'h000;
			{9'd134, 8'd127}: color_data = 12'h068;
			{9'd134, 8'd128}: color_data = 12'h079;
			{9'd134, 8'd129}: color_data = 12'h000;
			{9'd134, 8'd222}: color_data = 12'h200;
			{9'd134, 8'd223}: color_data = 12'h800;
			{9'd134, 8'd224}: color_data = 12'ha00;
			{9'd134, 8'd225}: color_data = 12'h700;
			{9'd134, 8'd226}: color_data = 12'h200;
			{9'd134, 8'd227}: color_data = 12'h920;
			{9'd134, 8'd228}: color_data = 12'hd30;
			{9'd134, 8'd229}: color_data = 12'h910;
			{9'd134, 8'd230}: color_data = 12'h200;
			{9'd134, 8'd231}: color_data = 12'h400;
			{9'd134, 8'd232}: color_data = 12'h900;
			{9'd134, 8'd233}: color_data = 12'ha00;
			{9'd134, 8'd234}: color_data = 12'h400;
			{9'd134, 8'd235}: color_data = 12'h310;
			{9'd134, 8'd236}: color_data = 12'hc30;
			{9'd134, 8'd237}: color_data = 12'hc20;
			{9'd134, 8'd238}: color_data = 12'h600;
			{9'd134, 8'd239}: color_data = 12'h000;
			{9'd135, 8'd68}: color_data = 12'h047;
			{9'd135, 8'd69}: color_data = 12'h6df;
			{9'd135, 8'd70}: color_data = 12'hfff;
			{9'd135, 8'd71}: color_data = 12'hcbb;
			{9'd135, 8'd72}: color_data = 12'h323;
			{9'd135, 8'd73}: color_data = 12'h002;
			{9'd135, 8'd74}: color_data = 12'h000;
			{9'd135, 8'd75}: color_data = 12'h012;
			{9'd135, 8'd76}: color_data = 12'h08c;
			{9'd135, 8'd77}: color_data = 12'h034;
			{9'd135, 8'd119}: color_data = 12'h000;
			{9'd135, 8'd120}: color_data = 12'h1ac;
			{9'd135, 8'd121}: color_data = 12'hdff;
			{9'd135, 8'd122}: color_data = 12'hfee;
			{9'd135, 8'd123}: color_data = 12'h666;
			{9'd135, 8'd124}: color_data = 12'h002;
			{9'd135, 8'd125}: color_data = 12'h001;
			{9'd135, 8'd126}: color_data = 12'h000;
			{9'd135, 8'd127}: color_data = 12'h068;
			{9'd135, 8'd128}: color_data = 12'h079;
			{9'd135, 8'd129}: color_data = 12'h000;
			{9'd135, 8'd222}: color_data = 12'h200;
			{9'd135, 8'd223}: color_data = 12'h900;
			{9'd135, 8'd224}: color_data = 12'ha00;
			{9'd135, 8'd225}: color_data = 12'h800;
			{9'd135, 8'd226}: color_data = 12'h100;
			{9'd135, 8'd227}: color_data = 12'h100;
			{9'd135, 8'd228}: color_data = 12'h300;
			{9'd135, 8'd229}: color_data = 12'h200;
			{9'd135, 8'd230}: color_data = 12'h000;
			{9'd135, 8'd231}: color_data = 12'h500;
			{9'd135, 8'd232}: color_data = 12'ha00;
			{9'd135, 8'd233}: color_data = 12'ha00;
			{9'd135, 8'd234}: color_data = 12'h500;
			{9'd135, 8'd235}: color_data = 12'h000;
			{9'd135, 8'd236}: color_data = 12'h200;
			{9'd135, 8'd237}: color_data = 12'h300;
			{9'd135, 8'd238}: color_data = 12'h100;
			{9'd135, 8'd239}: color_data = 12'h000;
			{9'd136, 8'd68}: color_data = 12'h047;
			{9'd136, 8'd69}: color_data = 12'h6ef;
			{9'd136, 8'd70}: color_data = 12'hddc;
			{9'd136, 8'd71}: color_data = 12'h434;
			{9'd136, 8'd72}: color_data = 12'h003;
			{9'd136, 8'd73}: color_data = 12'h005;
			{9'd136, 8'd74}: color_data = 12'h002;
			{9'd136, 8'd75}: color_data = 12'h012;
			{9'd136, 8'd76}: color_data = 12'h08c;
			{9'd136, 8'd77}: color_data = 12'h034;
			{9'd136, 8'd119}: color_data = 12'h000;
			{9'd136, 8'd120}: color_data = 12'h2ad;
			{9'd136, 8'd121}: color_data = 12'hcff;
			{9'd136, 8'd122}: color_data = 12'h877;
			{9'd136, 8'd123}: color_data = 12'h002;
			{9'd136, 8'd124}: color_data = 12'h004;
			{9'd136, 8'd125}: color_data = 12'h004;
			{9'd136, 8'd126}: color_data = 12'h000;
			{9'd136, 8'd127}: color_data = 12'h068;
			{9'd136, 8'd128}: color_data = 12'h079;
			{9'd136, 8'd129}: color_data = 12'h000;
			{9'd136, 8'd222}: color_data = 12'h300;
			{9'd136, 8'd223}: color_data = 12'hc20;
			{9'd136, 8'd224}: color_data = 12'ha00;
			{9'd136, 8'd225}: color_data = 12'h800;
			{9'd136, 8'd226}: color_data = 12'h100;
			{9'd136, 8'd227}: color_data = 12'h300;
			{9'd136, 8'd228}: color_data = 12'h500;
			{9'd136, 8'd229}: color_data = 12'h500;
			{9'd136, 8'd230}: color_data = 12'h100;
			{9'd136, 8'd231}: color_data = 12'h710;
			{9'd136, 8'd232}: color_data = 12'hc10;
			{9'd136, 8'd233}: color_data = 12'h900;
			{9'd136, 8'd234}: color_data = 12'h500;
			{9'd136, 8'd235}: color_data = 12'h100;
			{9'd136, 8'd236}: color_data = 12'h500;
			{9'd136, 8'd237}: color_data = 12'h600;
			{9'd136, 8'd238}: color_data = 12'h400;
			{9'd136, 8'd239}: color_data = 12'h000;
			{9'd137, 8'd68}: color_data = 12'h057;
			{9'd137, 8'd69}: color_data = 12'h3bd;
			{9'd137, 8'd70}: color_data = 12'h555;
			{9'd137, 8'd71}: color_data = 12'h002;
			{9'd137, 8'd72}: color_data = 12'h005;
			{9'd137, 8'd73}: color_data = 12'h005;
			{9'd137, 8'd74}: color_data = 12'h004;
			{9'd137, 8'd75}: color_data = 12'h025;
			{9'd137, 8'd76}: color_data = 12'h09c;
			{9'd137, 8'd77}: color_data = 12'h034;
			{9'd137, 8'd119}: color_data = 12'h000;
			{9'd137, 8'd120}: color_data = 12'h1ac;
			{9'd137, 8'd121}: color_data = 12'h689;
			{9'd137, 8'd122}: color_data = 12'h212;
			{9'd137, 8'd123}: color_data = 12'h004;
			{9'd137, 8'd124}: color_data = 12'h005;
			{9'd137, 8'd125}: color_data = 12'h005;
			{9'd137, 8'd126}: color_data = 12'h003;
			{9'd137, 8'd127}: color_data = 12'h06a;
			{9'd137, 8'd128}: color_data = 12'h079;
			{9'd137, 8'd129}: color_data = 12'h000;
			{9'd137, 8'd222}: color_data = 12'h410;
			{9'd137, 8'd223}: color_data = 12'hd30;
			{9'd137, 8'd224}: color_data = 12'hb00;
			{9'd137, 8'd225}: color_data = 12'h700;
			{9'd137, 8'd226}: color_data = 12'h200;
			{9'd137, 8'd227}: color_data = 12'h700;
			{9'd137, 8'd228}: color_data = 12'hb00;
			{9'd137, 8'd229}: color_data = 12'ha00;
			{9'd137, 8'd230}: color_data = 12'h300;
			{9'd137, 8'd231}: color_data = 12'h820;
			{9'd137, 8'd232}: color_data = 12'hd20;
			{9'd137, 8'd233}: color_data = 12'h900;
			{9'd137, 8'd234}: color_data = 12'h500;
			{9'd137, 8'd235}: color_data = 12'h300;
			{9'd137, 8'd236}: color_data = 12'h900;
			{9'd137, 8'd237}: color_data = 12'hb00;
			{9'd137, 8'd238}: color_data = 12'h800;
			{9'd137, 8'd239}: color_data = 12'h100;
			{9'd138, 8'd68}: color_data = 12'h046;
			{9'd138, 8'd69}: color_data = 12'h058;
			{9'd138, 8'd70}: color_data = 12'h002;
			{9'd138, 8'd71}: color_data = 12'h005;
			{9'd138, 8'd72}: color_data = 12'h005;
			{9'd138, 8'd73}: color_data = 12'h005;
			{9'd138, 8'd74}: color_data = 12'h005;
			{9'd138, 8'd75}: color_data = 12'h017;
			{9'd138, 8'd76}: color_data = 12'h05a;
			{9'd138, 8'd77}: color_data = 12'h023;
			{9'd138, 8'd119}: color_data = 12'h000;
			{9'd138, 8'd120}: color_data = 12'h058;
			{9'd138, 8'd121}: color_data = 12'h013;
			{9'd138, 8'd122}: color_data = 12'h002;
			{9'd138, 8'd123}: color_data = 12'h004;
			{9'd138, 8'd124}: color_data = 12'h004;
			{9'd138, 8'd125}: color_data = 12'h004;
			{9'd138, 8'd126}: color_data = 12'h004;
			{9'd138, 8'd127}: color_data = 12'h039;
			{9'd138, 8'd128}: color_data = 12'h046;
			{9'd138, 8'd129}: color_data = 12'h000;
			{9'd138, 8'd222}: color_data = 12'h410;
			{9'd138, 8'd223}: color_data = 12'he40;
			{9'd138, 8'd224}: color_data = 12'hd20;
			{9'd138, 8'd225}: color_data = 12'h800;
			{9'd138, 8'd226}: color_data = 12'h200;
			{9'd138, 8'd227}: color_data = 12'h600;
			{9'd138, 8'd228}: color_data = 12'ha00;
			{9'd138, 8'd229}: color_data = 12'h900;
			{9'd138, 8'd230}: color_data = 12'h300;
			{9'd138, 8'd231}: color_data = 12'h820;
			{9'd138, 8'd232}: color_data = 12'hf30;
			{9'd138, 8'd233}: color_data = 12'hc00;
			{9'd138, 8'd234}: color_data = 12'h500;
			{9'd138, 8'd235}: color_data = 12'h200;
			{9'd138, 8'd236}: color_data = 12'h900;
			{9'd138, 8'd237}: color_data = 12'ha00;
			{9'd138, 8'd238}: color_data = 12'h700;
			{9'd138, 8'd239}: color_data = 12'h100;
			{9'd139, 8'd68}: color_data = 12'h002;
			{9'd139, 8'd69}: color_data = 12'h004;
			{9'd139, 8'd70}: color_data = 12'h004;
			{9'd139, 8'd71}: color_data = 12'h004;
			{9'd139, 8'd72}: color_data = 12'h004;
			{9'd139, 8'd73}: color_data = 12'h004;
			{9'd139, 8'd74}: color_data = 12'h004;
			{9'd139, 8'd75}: color_data = 12'h004;
			{9'd139, 8'd76}: color_data = 12'h004;
			{9'd139, 8'd77}: color_data = 12'h001;
			{9'd139, 8'd119}: color_data = 12'h000;
			{9'd139, 8'd120}: color_data = 12'h016;
			{9'd139, 8'd121}: color_data = 12'h017;
			{9'd139, 8'd122}: color_data = 12'h017;
			{9'd139, 8'd123}: color_data = 12'h027;
			{9'd139, 8'd124}: color_data = 12'h027;
			{9'd139, 8'd125}: color_data = 12'h027;
			{9'd139, 8'd126}: color_data = 12'h027;
			{9'd139, 8'd127}: color_data = 12'h028;
			{9'd139, 8'd128}: color_data = 12'h014;
			{9'd139, 8'd129}: color_data = 12'h000;
			{9'd139, 8'd222}: color_data = 12'h300;
			{9'd139, 8'd223}: color_data = 12'hc30;
			{9'd139, 8'd224}: color_data = 12'hc30;
			{9'd139, 8'd225}: color_data = 12'h600;
			{9'd139, 8'd226}: color_data = 12'h100;
			{9'd139, 8'd227}: color_data = 12'h600;
			{9'd139, 8'd228}: color_data = 12'ha00;
			{9'd139, 8'd229}: color_data = 12'h900;
			{9'd139, 8'd230}: color_data = 12'h300;
			{9'd139, 8'd231}: color_data = 12'h620;
			{9'd139, 8'd232}: color_data = 12'hd40;
			{9'd139, 8'd233}: color_data = 12'ha20;
			{9'd139, 8'd234}: color_data = 12'h300;
			{9'd139, 8'd235}: color_data = 12'h200;
			{9'd139, 8'd236}: color_data = 12'h900;
			{9'd139, 8'd237}: color_data = 12'ha00;
			{9'd139, 8'd238}: color_data = 12'h700;
			{9'd139, 8'd239}: color_data = 12'h100;
			{9'd140, 8'd68}: color_data = 12'h000;
			{9'd140, 8'd69}: color_data = 12'h000;
			{9'd140, 8'd70}: color_data = 12'h001;
			{9'd140, 8'd71}: color_data = 12'h000;
			{9'd140, 8'd72}: color_data = 12'h000;
			{9'd140, 8'd73}: color_data = 12'h000;
			{9'd140, 8'd74}: color_data = 12'h000;
			{9'd140, 8'd75}: color_data = 12'h000;
			{9'd140, 8'd76}: color_data = 12'h000;
			{9'd140, 8'd77}: color_data = 12'h000;
			{9'd140, 8'd119}: color_data = 12'h000;
			{9'd140, 8'd120}: color_data = 12'h07b;
			{9'd140, 8'd121}: color_data = 12'h0ae;
			{9'd140, 8'd122}: color_data = 12'h09e;
			{9'd140, 8'd123}: color_data = 12'h09e;
			{9'd140, 8'd124}: color_data = 12'h09e;
			{9'd140, 8'd125}: color_data = 12'h09e;
			{9'd140, 8'd126}: color_data = 12'h09e;
			{9'd140, 8'd127}: color_data = 12'h09e;
			{9'd140, 8'd128}: color_data = 12'h057;
			{9'd140, 8'd129}: color_data = 12'h000;
			{9'd140, 8'd222}: color_data = 12'h000;
			{9'd140, 8'd223}: color_data = 12'h200;
			{9'd140, 8'd224}: color_data = 12'h300;
			{9'd140, 8'd225}: color_data = 12'h100;
			{9'd140, 8'd226}: color_data = 12'h000;
			{9'd140, 8'd227}: color_data = 12'h700;
			{9'd140, 8'd228}: color_data = 12'ha00;
			{9'd140, 8'd229}: color_data = 12'h900;
			{9'd140, 8'd230}: color_data = 12'h300;
			{9'd140, 8'd231}: color_data = 12'h100;
			{9'd140, 8'd232}: color_data = 12'h310;
			{9'd140, 8'd233}: color_data = 12'h200;
			{9'd140, 8'd234}: color_data = 12'h000;
			{9'd140, 8'd235}: color_data = 12'h300;
			{9'd140, 8'd236}: color_data = 12'h900;
			{9'd140, 8'd237}: color_data = 12'ha00;
			{9'd140, 8'd238}: color_data = 12'h700;
			{9'd140, 8'd239}: color_data = 12'h100;
			{9'd141, 8'd119}: color_data = 12'h000;
			{9'd141, 8'd120}: color_data = 12'h1ad;
			{9'd141, 8'd121}: color_data = 12'h8ff;
			{9'd141, 8'd122}: color_data = 12'h3df;
			{9'd141, 8'd123}: color_data = 12'h0bf;
			{9'd141, 8'd124}: color_data = 12'h0cf;
			{9'd141, 8'd125}: color_data = 12'h0cf;
			{9'd141, 8'd126}: color_data = 12'h07a;
			{9'd141, 8'd127}: color_data = 12'h08b;
			{9'd141, 8'd128}: color_data = 12'h079;
			{9'd141, 8'd129}: color_data = 12'h000;
			{9'd141, 8'd222}: color_data = 12'h100;
			{9'd141, 8'd223}: color_data = 12'h400;
			{9'd141, 8'd224}: color_data = 12'h500;
			{9'd141, 8'd225}: color_data = 12'h400;
			{9'd141, 8'd226}: color_data = 12'h200;
			{9'd141, 8'd227}: color_data = 12'ha20;
			{9'd141, 8'd228}: color_data = 12'hb10;
			{9'd141, 8'd229}: color_data = 12'h900;
			{9'd141, 8'd230}: color_data = 12'h300;
			{9'd141, 8'd231}: color_data = 12'h200;
			{9'd141, 8'd232}: color_data = 12'h500;
			{9'd141, 8'd233}: color_data = 12'h500;
			{9'd141, 8'd234}: color_data = 12'h200;
			{9'd141, 8'd235}: color_data = 12'h410;
			{9'd141, 8'd236}: color_data = 12'hc20;
			{9'd141, 8'd237}: color_data = 12'ha00;
			{9'd141, 8'd238}: color_data = 12'h700;
			{9'd141, 8'd239}: color_data = 12'h100;
			{9'd142, 8'd119}: color_data = 12'h000;
			{9'd142, 8'd120}: color_data = 12'h2ac;
			{9'd142, 8'd121}: color_data = 12'hdff;
			{9'd142, 8'd122}: color_data = 12'haef;
			{9'd142, 8'd123}: color_data = 12'h1bf;
			{9'd142, 8'd124}: color_data = 12'h0cf;
			{9'd142, 8'd125}: color_data = 12'h08b;
			{9'd142, 8'd126}: color_data = 12'h012;
			{9'd142, 8'd127}: color_data = 12'h068;
			{9'd142, 8'd128}: color_data = 12'h079;
			{9'd142, 8'd129}: color_data = 12'h000;
			{9'd142, 8'd222}: color_data = 12'h200;
			{9'd142, 8'd223}: color_data = 12'h900;
			{9'd142, 8'd224}: color_data = 12'hb00;
			{9'd142, 8'd225}: color_data = 12'h800;
			{9'd142, 8'd226}: color_data = 12'h200;
			{9'd142, 8'd227}: color_data = 12'hb30;
			{9'd142, 8'd228}: color_data = 12'hc10;
			{9'd142, 8'd229}: color_data = 12'h800;
			{9'd142, 8'd230}: color_data = 12'h300;
			{9'd142, 8'd231}: color_data = 12'h400;
			{9'd142, 8'd232}: color_data = 12'ha00;
			{9'd142, 8'd233}: color_data = 12'ha00;
			{9'd142, 8'd234}: color_data = 12'h500;
			{9'd142, 8'd235}: color_data = 12'h510;
			{9'd142, 8'd236}: color_data = 12'hd30;
			{9'd142, 8'd237}: color_data = 12'ha00;
			{9'd142, 8'd238}: color_data = 12'h700;
			{9'd142, 8'd239}: color_data = 12'h100;
			{9'd143, 8'd119}: color_data = 12'h000;
			{9'd143, 8'd120}: color_data = 12'h1ac;
			{9'd143, 8'd121}: color_data = 12'hdff;
			{9'd143, 8'd122}: color_data = 12'hfff;
			{9'd143, 8'd123}: color_data = 12'h8ef;
			{9'd143, 8'd124}: color_data = 12'h19c;
			{9'd143, 8'd125}: color_data = 12'h023;
			{9'd143, 8'd127}: color_data = 12'h068;
			{9'd143, 8'd128}: color_data = 12'h079;
			{9'd143, 8'd129}: color_data = 12'h000;
			{9'd143, 8'd222}: color_data = 12'h200;
			{9'd143, 8'd223}: color_data = 12'h900;
			{9'd143, 8'd224}: color_data = 12'ha00;
			{9'd143, 8'd225}: color_data = 12'h700;
			{9'd143, 8'd226}: color_data = 12'h200;
			{9'd143, 8'd227}: color_data = 12'hb30;
			{9'd143, 8'd228}: color_data = 12'he20;
			{9'd143, 8'd229}: color_data = 12'ha00;
			{9'd143, 8'd230}: color_data = 12'h300;
			{9'd143, 8'd231}: color_data = 12'h400;
			{9'd143, 8'd232}: color_data = 12'ha00;
			{9'd143, 8'd233}: color_data = 12'ha00;
			{9'd143, 8'd234}: color_data = 12'h400;
			{9'd143, 8'd235}: color_data = 12'h510;
			{9'd143, 8'd236}: color_data = 12'hf40;
			{9'd143, 8'd237}: color_data = 12'hd10;
			{9'd143, 8'd238}: color_data = 12'h800;
			{9'd143, 8'd239}: color_data = 12'h100;
			{9'd144, 8'd119}: color_data = 12'h000;
			{9'd144, 8'd120}: color_data = 12'h1ac;
			{9'd144, 8'd121}: color_data = 12'hcff;
			{9'd144, 8'd122}: color_data = 12'hfff;
			{9'd144, 8'd123}: color_data = 12'hddd;
			{9'd144, 8'd124}: color_data = 12'h345;
			{9'd144, 8'd126}: color_data = 12'h000;
			{9'd144, 8'd127}: color_data = 12'h068;
			{9'd144, 8'd128}: color_data = 12'h079;
			{9'd144, 8'd129}: color_data = 12'h000;
			{9'd144, 8'd222}: color_data = 12'h200;
			{9'd144, 8'd223}: color_data = 12'h800;
			{9'd144, 8'd224}: color_data = 12'ha00;
			{9'd144, 8'd225}: color_data = 12'h700;
			{9'd144, 8'd226}: color_data = 12'h200;
			{9'd144, 8'd227}: color_data = 12'h920;
			{9'd144, 8'd228}: color_data = 12'hd30;
			{9'd144, 8'd229}: color_data = 12'h910;
			{9'd144, 8'd230}: color_data = 12'h200;
			{9'd144, 8'd231}: color_data = 12'h400;
			{9'd144, 8'd232}: color_data = 12'h900;
			{9'd144, 8'd233}: color_data = 12'ha00;
			{9'd144, 8'd234}: color_data = 12'h400;
			{9'd144, 8'd235}: color_data = 12'h310;
			{9'd144, 8'd236}: color_data = 12'hc30;
			{9'd144, 8'd237}: color_data = 12'hc20;
			{9'd144, 8'd238}: color_data = 12'h600;
			{9'd144, 8'd239}: color_data = 12'h000;
			{9'd145, 8'd119}: color_data = 12'h000;
			{9'd145, 8'd120}: color_data = 12'h1ac;
			{9'd145, 8'd121}: color_data = 12'hdff;
			{9'd145, 8'd122}: color_data = 12'hfee;
			{9'd145, 8'd123}: color_data = 12'h666;
			{9'd145, 8'd124}: color_data = 12'h002;
			{9'd145, 8'd125}: color_data = 12'h001;
			{9'd145, 8'd126}: color_data = 12'h000;
			{9'd145, 8'd127}: color_data = 12'h068;
			{9'd145, 8'd128}: color_data = 12'h079;
			{9'd145, 8'd129}: color_data = 12'h000;
			{9'd145, 8'd222}: color_data = 12'h200;
			{9'd145, 8'd223}: color_data = 12'h900;
			{9'd145, 8'd224}: color_data = 12'ha00;
			{9'd145, 8'd225}: color_data = 12'h800;
			{9'd145, 8'd226}: color_data = 12'h100;
			{9'd145, 8'd227}: color_data = 12'h100;
			{9'd145, 8'd228}: color_data = 12'h310;
			{9'd145, 8'd229}: color_data = 12'h200;
			{9'd145, 8'd230}: color_data = 12'h000;
			{9'd145, 8'd231}: color_data = 12'h500;
			{9'd145, 8'd232}: color_data = 12'ha00;
			{9'd145, 8'd233}: color_data = 12'ha00;
			{9'd145, 8'd234}: color_data = 12'h500;
			{9'd145, 8'd235}: color_data = 12'h000;
			{9'd145, 8'd236}: color_data = 12'h200;
			{9'd145, 8'd237}: color_data = 12'h300;
			{9'd145, 8'd238}: color_data = 12'h100;
			{9'd145, 8'd239}: color_data = 12'h000;
			{9'd146, 8'd119}: color_data = 12'h000;
			{9'd146, 8'd120}: color_data = 12'h2ad;
			{9'd146, 8'd121}: color_data = 12'hcff;
			{9'd146, 8'd122}: color_data = 12'h877;
			{9'd146, 8'd123}: color_data = 12'h002;
			{9'd146, 8'd124}: color_data = 12'h004;
			{9'd146, 8'd125}: color_data = 12'h004;
			{9'd146, 8'd126}: color_data = 12'h000;
			{9'd146, 8'd127}: color_data = 12'h068;
			{9'd146, 8'd128}: color_data = 12'h079;
			{9'd146, 8'd129}: color_data = 12'h000;
			{9'd146, 8'd222}: color_data = 12'h300;
			{9'd146, 8'd223}: color_data = 12'hc20;
			{9'd146, 8'd224}: color_data = 12'ha00;
			{9'd146, 8'd225}: color_data = 12'h800;
			{9'd146, 8'd226}: color_data = 12'h100;
			{9'd146, 8'd227}: color_data = 12'h300;
			{9'd146, 8'd228}: color_data = 12'h500;
			{9'd146, 8'd229}: color_data = 12'h500;
			{9'd146, 8'd230}: color_data = 12'h100;
			{9'd146, 8'd231}: color_data = 12'h710;
			{9'd146, 8'd232}: color_data = 12'hc10;
			{9'd146, 8'd233}: color_data = 12'h900;
			{9'd146, 8'd234}: color_data = 12'h500;
			{9'd146, 8'd235}: color_data = 12'h100;
			{9'd146, 8'd236}: color_data = 12'h500;
			{9'd146, 8'd237}: color_data = 12'h600;
			{9'd146, 8'd238}: color_data = 12'h400;
			{9'd146, 8'd239}: color_data = 12'h000;
			{9'd147, 8'd119}: color_data = 12'h000;
			{9'd147, 8'd120}: color_data = 12'h1ac;
			{9'd147, 8'd121}: color_data = 12'h689;
			{9'd147, 8'd122}: color_data = 12'h212;
			{9'd147, 8'd123}: color_data = 12'h004;
			{9'd147, 8'd124}: color_data = 12'h005;
			{9'd147, 8'd125}: color_data = 12'h005;
			{9'd147, 8'd126}: color_data = 12'h003;
			{9'd147, 8'd127}: color_data = 12'h06a;
			{9'd147, 8'd128}: color_data = 12'h079;
			{9'd147, 8'd129}: color_data = 12'h000;
			{9'd147, 8'd222}: color_data = 12'h410;
			{9'd147, 8'd223}: color_data = 12'hd30;
			{9'd147, 8'd224}: color_data = 12'hb00;
			{9'd147, 8'd225}: color_data = 12'h700;
			{9'd147, 8'd226}: color_data = 12'h200;
			{9'd147, 8'd227}: color_data = 12'h700;
			{9'd147, 8'd228}: color_data = 12'hb00;
			{9'd147, 8'd229}: color_data = 12'ha00;
			{9'd147, 8'd230}: color_data = 12'h300;
			{9'd147, 8'd231}: color_data = 12'h820;
			{9'd147, 8'd232}: color_data = 12'hd20;
			{9'd147, 8'd233}: color_data = 12'h900;
			{9'd147, 8'd234}: color_data = 12'h500;
			{9'd147, 8'd235}: color_data = 12'h300;
			{9'd147, 8'd236}: color_data = 12'h900;
			{9'd147, 8'd237}: color_data = 12'hb00;
			{9'd147, 8'd238}: color_data = 12'h800;
			{9'd147, 8'd239}: color_data = 12'h100;
			{9'd148, 8'd119}: color_data = 12'h000;
			{9'd148, 8'd120}: color_data = 12'h058;
			{9'd148, 8'd121}: color_data = 12'h013;
			{9'd148, 8'd122}: color_data = 12'h002;
			{9'd148, 8'd123}: color_data = 12'h004;
			{9'd148, 8'd124}: color_data = 12'h004;
			{9'd148, 8'd125}: color_data = 12'h004;
			{9'd148, 8'd126}: color_data = 12'h004;
			{9'd148, 8'd127}: color_data = 12'h039;
			{9'd148, 8'd128}: color_data = 12'h046;
			{9'd148, 8'd129}: color_data = 12'h000;
			{9'd148, 8'd222}: color_data = 12'h410;
			{9'd148, 8'd223}: color_data = 12'he40;
			{9'd148, 8'd224}: color_data = 12'hd20;
			{9'd148, 8'd225}: color_data = 12'h800;
			{9'd148, 8'd226}: color_data = 12'h200;
			{9'd148, 8'd227}: color_data = 12'h600;
			{9'd148, 8'd228}: color_data = 12'ha00;
			{9'd148, 8'd229}: color_data = 12'h900;
			{9'd148, 8'd230}: color_data = 12'h300;
			{9'd148, 8'd231}: color_data = 12'h820;
			{9'd148, 8'd232}: color_data = 12'hf30;
			{9'd148, 8'd233}: color_data = 12'hc00;
			{9'd148, 8'd234}: color_data = 12'h500;
			{9'd148, 8'd235}: color_data = 12'h200;
			{9'd148, 8'd236}: color_data = 12'h900;
			{9'd148, 8'd237}: color_data = 12'ha00;
			{9'd148, 8'd238}: color_data = 12'h700;
			{9'd148, 8'd239}: color_data = 12'h100;
			{9'd149, 8'd119}: color_data = 12'h000;
			{9'd149, 8'd120}: color_data = 12'h016;
			{9'd149, 8'd121}: color_data = 12'h017;
			{9'd149, 8'd122}: color_data = 12'h016;
			{9'd149, 8'd123}: color_data = 12'h027;
			{9'd149, 8'd124}: color_data = 12'h027;
			{9'd149, 8'd125}: color_data = 12'h027;
			{9'd149, 8'd126}: color_data = 12'h027;
			{9'd149, 8'd127}: color_data = 12'h028;
			{9'd149, 8'd128}: color_data = 12'h014;
			{9'd149, 8'd129}: color_data = 12'h000;
			{9'd149, 8'd222}: color_data = 12'h300;
			{9'd149, 8'd223}: color_data = 12'hc30;
			{9'd149, 8'd224}: color_data = 12'hc30;
			{9'd149, 8'd225}: color_data = 12'h700;
			{9'd149, 8'd226}: color_data = 12'h100;
			{9'd149, 8'd227}: color_data = 12'h600;
			{9'd149, 8'd228}: color_data = 12'ha00;
			{9'd149, 8'd229}: color_data = 12'h900;
			{9'd149, 8'd230}: color_data = 12'h300;
			{9'd149, 8'd231}: color_data = 12'h620;
			{9'd149, 8'd232}: color_data = 12'hd40;
			{9'd149, 8'd233}: color_data = 12'ha20;
			{9'd149, 8'd234}: color_data = 12'h300;
			{9'd149, 8'd235}: color_data = 12'h200;
			{9'd149, 8'd236}: color_data = 12'h800;
			{9'd149, 8'd237}: color_data = 12'ha00;
			{9'd149, 8'd238}: color_data = 12'h700;
			{9'd149, 8'd239}: color_data = 12'h100;
			{9'd150, 8'd119}: color_data = 12'h000;
			{9'd150, 8'd120}: color_data = 12'h07b;
			{9'd150, 8'd121}: color_data = 12'h0ae;
			{9'd150, 8'd122}: color_data = 12'h09e;
			{9'd150, 8'd123}: color_data = 12'h09e;
			{9'd150, 8'd124}: color_data = 12'h09e;
			{9'd150, 8'd125}: color_data = 12'h09e;
			{9'd150, 8'd126}: color_data = 12'h09e;
			{9'd150, 8'd127}: color_data = 12'h09e;
			{9'd150, 8'd128}: color_data = 12'h057;
			{9'd150, 8'd129}: color_data = 12'h000;
			{9'd150, 8'd222}: color_data = 12'h000;
			{9'd150, 8'd223}: color_data = 12'h200;
			{9'd150, 8'd224}: color_data = 12'h300;
			{9'd150, 8'd225}: color_data = 12'h100;
			{9'd150, 8'd226}: color_data = 12'h000;
			{9'd150, 8'd227}: color_data = 12'h700;
			{9'd150, 8'd228}: color_data = 12'ha00;
			{9'd150, 8'd229}: color_data = 12'h900;
			{9'd150, 8'd230}: color_data = 12'h300;
			{9'd150, 8'd231}: color_data = 12'h100;
			{9'd150, 8'd232}: color_data = 12'h310;
			{9'd150, 8'd233}: color_data = 12'h200;
			{9'd150, 8'd234}: color_data = 12'h000;
			{9'd150, 8'd235}: color_data = 12'h300;
			{9'd150, 8'd236}: color_data = 12'h900;
			{9'd150, 8'd237}: color_data = 12'ha00;
			{9'd150, 8'd238}: color_data = 12'h700;
			{9'd150, 8'd239}: color_data = 12'h100;
			{9'd151, 8'd119}: color_data = 12'h000;
			{9'd151, 8'd120}: color_data = 12'h1ad;
			{9'd151, 8'd121}: color_data = 12'h8ff;
			{9'd151, 8'd122}: color_data = 12'h3df;
			{9'd151, 8'd123}: color_data = 12'h0cf;
			{9'd151, 8'd124}: color_data = 12'h0cf;
			{9'd151, 8'd125}: color_data = 12'h0cf;
			{9'd151, 8'd126}: color_data = 12'h079;
			{9'd151, 8'd127}: color_data = 12'h08b;
			{9'd151, 8'd128}: color_data = 12'h079;
			{9'd151, 8'd129}: color_data = 12'h000;
			{9'd151, 8'd222}: color_data = 12'h100;
			{9'd151, 8'd223}: color_data = 12'h500;
			{9'd151, 8'd224}: color_data = 12'h500;
			{9'd151, 8'd225}: color_data = 12'h400;
			{9'd151, 8'd226}: color_data = 12'h100;
			{9'd151, 8'd227}: color_data = 12'ha20;
			{9'd151, 8'd228}: color_data = 12'hb10;
			{9'd151, 8'd229}: color_data = 12'h900;
			{9'd151, 8'd230}: color_data = 12'h300;
			{9'd151, 8'd231}: color_data = 12'h200;
			{9'd151, 8'd232}: color_data = 12'h500;
			{9'd151, 8'd233}: color_data = 12'h500;
			{9'd151, 8'd234}: color_data = 12'h200;
			{9'd151, 8'd235}: color_data = 12'h410;
			{9'd151, 8'd236}: color_data = 12'hc20;
			{9'd151, 8'd237}: color_data = 12'ha00;
			{9'd151, 8'd238}: color_data = 12'h700;
			{9'd151, 8'd239}: color_data = 12'h100;
			{9'd152, 8'd119}: color_data = 12'h000;
			{9'd152, 8'd120}: color_data = 12'h2ac;
			{9'd152, 8'd121}: color_data = 12'hdff;
			{9'd152, 8'd122}: color_data = 12'haef;
			{9'd152, 8'd123}: color_data = 12'h1cf;
			{9'd152, 8'd124}: color_data = 12'h0cf;
			{9'd152, 8'd125}: color_data = 12'h08b;
			{9'd152, 8'd126}: color_data = 12'h012;
			{9'd152, 8'd127}: color_data = 12'h068;
			{9'd152, 8'd128}: color_data = 12'h079;
			{9'd152, 8'd129}: color_data = 12'h000;
			{9'd152, 8'd222}: color_data = 12'h200;
			{9'd152, 8'd223}: color_data = 12'h900;
			{9'd152, 8'd224}: color_data = 12'hb00;
			{9'd152, 8'd225}: color_data = 12'h800;
			{9'd152, 8'd226}: color_data = 12'h200;
			{9'd152, 8'd227}: color_data = 12'hb30;
			{9'd152, 8'd228}: color_data = 12'hc10;
			{9'd152, 8'd229}: color_data = 12'h800;
			{9'd152, 8'd230}: color_data = 12'h300;
			{9'd152, 8'd231}: color_data = 12'h400;
			{9'd152, 8'd232}: color_data = 12'ha00;
			{9'd152, 8'd233}: color_data = 12'ha00;
			{9'd152, 8'd234}: color_data = 12'h500;
			{9'd152, 8'd235}: color_data = 12'h510;
			{9'd152, 8'd236}: color_data = 12'hd30;
			{9'd152, 8'd237}: color_data = 12'ha00;
			{9'd152, 8'd238}: color_data = 12'h700;
			{9'd152, 8'd239}: color_data = 12'h100;
			{9'd153, 8'd119}: color_data = 12'h000;
			{9'd153, 8'd120}: color_data = 12'h1ac;
			{9'd153, 8'd121}: color_data = 12'hdff;
			{9'd153, 8'd122}: color_data = 12'hfff;
			{9'd153, 8'd123}: color_data = 12'h8ef;
			{9'd153, 8'd124}: color_data = 12'h19c;
			{9'd153, 8'd125}: color_data = 12'h023;
			{9'd153, 8'd127}: color_data = 12'h068;
			{9'd153, 8'd128}: color_data = 12'h079;
			{9'd153, 8'd129}: color_data = 12'h000;
			{9'd153, 8'd222}: color_data = 12'h200;
			{9'd153, 8'd223}: color_data = 12'h900;
			{9'd153, 8'd224}: color_data = 12'ha00;
			{9'd153, 8'd225}: color_data = 12'h700;
			{9'd153, 8'd226}: color_data = 12'h200;
			{9'd153, 8'd227}: color_data = 12'hb30;
			{9'd153, 8'd228}: color_data = 12'he20;
			{9'd153, 8'd229}: color_data = 12'ha00;
			{9'd153, 8'd230}: color_data = 12'h300;
			{9'd153, 8'd231}: color_data = 12'h400;
			{9'd153, 8'd232}: color_data = 12'ha00;
			{9'd153, 8'd233}: color_data = 12'ha00;
			{9'd153, 8'd234}: color_data = 12'h400;
			{9'd153, 8'd235}: color_data = 12'h510;
			{9'd153, 8'd236}: color_data = 12'hf40;
			{9'd153, 8'd237}: color_data = 12'hd10;
			{9'd153, 8'd238}: color_data = 12'h800;
			{9'd153, 8'd239}: color_data = 12'h100;
			{9'd154, 8'd119}: color_data = 12'h000;
			{9'd154, 8'd120}: color_data = 12'h1ac;
			{9'd154, 8'd121}: color_data = 12'hcff;
			{9'd154, 8'd122}: color_data = 12'hfff;
			{9'd154, 8'd123}: color_data = 12'hddd;
			{9'd154, 8'd124}: color_data = 12'h345;
			{9'd154, 8'd126}: color_data = 12'h000;
			{9'd154, 8'd127}: color_data = 12'h068;
			{9'd154, 8'd128}: color_data = 12'h079;
			{9'd154, 8'd129}: color_data = 12'h000;
			{9'd154, 8'd222}: color_data = 12'h200;
			{9'd154, 8'd223}: color_data = 12'h800;
			{9'd154, 8'd224}: color_data = 12'ha00;
			{9'd154, 8'd225}: color_data = 12'h800;
			{9'd154, 8'd226}: color_data = 12'h200;
			{9'd154, 8'd227}: color_data = 12'h920;
			{9'd154, 8'd228}: color_data = 12'hd30;
			{9'd154, 8'd229}: color_data = 12'h910;
			{9'd154, 8'd230}: color_data = 12'h200;
			{9'd154, 8'd231}: color_data = 12'h400;
			{9'd154, 8'd232}: color_data = 12'h900;
			{9'd154, 8'd233}: color_data = 12'ha00;
			{9'd154, 8'd234}: color_data = 12'h400;
			{9'd154, 8'd235}: color_data = 12'h310;
			{9'd154, 8'd236}: color_data = 12'hc30;
			{9'd154, 8'd237}: color_data = 12'hc20;
			{9'd154, 8'd238}: color_data = 12'h600;
			{9'd154, 8'd239}: color_data = 12'h000;
			{9'd155, 8'd119}: color_data = 12'h000;
			{9'd155, 8'd120}: color_data = 12'h1ac;
			{9'd155, 8'd121}: color_data = 12'hdff;
			{9'd155, 8'd122}: color_data = 12'hfee;
			{9'd155, 8'd123}: color_data = 12'h666;
			{9'd155, 8'd124}: color_data = 12'h002;
			{9'd155, 8'd125}: color_data = 12'h001;
			{9'd155, 8'd126}: color_data = 12'h000;
			{9'd155, 8'd127}: color_data = 12'h068;
			{9'd155, 8'd128}: color_data = 12'h079;
			{9'd155, 8'd129}: color_data = 12'h000;
			{9'd155, 8'd222}: color_data = 12'h200;
			{9'd155, 8'd223}: color_data = 12'h900;
			{9'd155, 8'd224}: color_data = 12'ha00;
			{9'd155, 8'd225}: color_data = 12'h800;
			{9'd155, 8'd226}: color_data = 12'h100;
			{9'd155, 8'd227}: color_data = 12'h100;
			{9'd155, 8'd228}: color_data = 12'h310;
			{9'd155, 8'd229}: color_data = 12'h200;
			{9'd155, 8'd230}: color_data = 12'h000;
			{9'd155, 8'd231}: color_data = 12'h500;
			{9'd155, 8'd232}: color_data = 12'ha00;
			{9'd155, 8'd233}: color_data = 12'ha00;
			{9'd155, 8'd234}: color_data = 12'h500;
			{9'd155, 8'd235}: color_data = 12'h000;
			{9'd155, 8'd236}: color_data = 12'h200;
			{9'd155, 8'd237}: color_data = 12'h300;
			{9'd155, 8'd238}: color_data = 12'h100;
			{9'd155, 8'd239}: color_data = 12'h000;
			{9'd156, 8'd119}: color_data = 12'h000;
			{9'd156, 8'd120}: color_data = 12'h2ad;
			{9'd156, 8'd121}: color_data = 12'hcff;
			{9'd156, 8'd122}: color_data = 12'h877;
			{9'd156, 8'd123}: color_data = 12'h002;
			{9'd156, 8'd124}: color_data = 12'h004;
			{9'd156, 8'd125}: color_data = 12'h004;
			{9'd156, 8'd126}: color_data = 12'h000;
			{9'd156, 8'd127}: color_data = 12'h068;
			{9'd156, 8'd128}: color_data = 12'h079;
			{9'd156, 8'd129}: color_data = 12'h000;
			{9'd156, 8'd222}: color_data = 12'h300;
			{9'd156, 8'd223}: color_data = 12'hc20;
			{9'd156, 8'd224}: color_data = 12'ha00;
			{9'd156, 8'd225}: color_data = 12'h800;
			{9'd156, 8'd226}: color_data = 12'h100;
			{9'd156, 8'd227}: color_data = 12'h300;
			{9'd156, 8'd228}: color_data = 12'h500;
			{9'd156, 8'd229}: color_data = 12'h500;
			{9'd156, 8'd230}: color_data = 12'h100;
			{9'd156, 8'd231}: color_data = 12'h710;
			{9'd156, 8'd232}: color_data = 12'hc10;
			{9'd156, 8'd233}: color_data = 12'h900;
			{9'd156, 8'd234}: color_data = 12'h500;
			{9'd156, 8'd235}: color_data = 12'h100;
			{9'd156, 8'd236}: color_data = 12'h500;
			{9'd156, 8'd237}: color_data = 12'h500;
			{9'd156, 8'd238}: color_data = 12'h400;
			{9'd156, 8'd239}: color_data = 12'h000;
			{9'd157, 8'd119}: color_data = 12'h000;
			{9'd157, 8'd120}: color_data = 12'h1ac;
			{9'd157, 8'd121}: color_data = 12'h689;
			{9'd157, 8'd122}: color_data = 12'h212;
			{9'd157, 8'd123}: color_data = 12'h004;
			{9'd157, 8'd124}: color_data = 12'h005;
			{9'd157, 8'd125}: color_data = 12'h005;
			{9'd157, 8'd126}: color_data = 12'h003;
			{9'd157, 8'd127}: color_data = 12'h06a;
			{9'd157, 8'd128}: color_data = 12'h079;
			{9'd157, 8'd129}: color_data = 12'h000;
			{9'd157, 8'd222}: color_data = 12'h410;
			{9'd157, 8'd223}: color_data = 12'hd30;
			{9'd157, 8'd224}: color_data = 12'hb00;
			{9'd157, 8'd225}: color_data = 12'h700;
			{9'd157, 8'd226}: color_data = 12'h200;
			{9'd157, 8'd227}: color_data = 12'h700;
			{9'd157, 8'd228}: color_data = 12'hb00;
			{9'd157, 8'd229}: color_data = 12'h900;
			{9'd157, 8'd230}: color_data = 12'h300;
			{9'd157, 8'd231}: color_data = 12'h820;
			{9'd157, 8'd232}: color_data = 12'hd20;
			{9'd157, 8'd233}: color_data = 12'h900;
			{9'd157, 8'd234}: color_data = 12'h500;
			{9'd157, 8'd235}: color_data = 12'h300;
			{9'd157, 8'd236}: color_data = 12'h900;
			{9'd157, 8'd237}: color_data = 12'hb00;
			{9'd157, 8'd238}: color_data = 12'h800;
			{9'd157, 8'd239}: color_data = 12'h100;
			{9'd158, 8'd119}: color_data = 12'h000;
			{9'd158, 8'd120}: color_data = 12'h058;
			{9'd158, 8'd121}: color_data = 12'h013;
			{9'd158, 8'd122}: color_data = 12'h002;
			{9'd158, 8'd123}: color_data = 12'h004;
			{9'd158, 8'd124}: color_data = 12'h004;
			{9'd158, 8'd125}: color_data = 12'h004;
			{9'd158, 8'd126}: color_data = 12'h004;
			{9'd158, 8'd127}: color_data = 12'h038;
			{9'd158, 8'd128}: color_data = 12'h046;
			{9'd158, 8'd129}: color_data = 12'h000;
			{9'd158, 8'd222}: color_data = 12'h410;
			{9'd158, 8'd223}: color_data = 12'he40;
			{9'd158, 8'd224}: color_data = 12'hd20;
			{9'd158, 8'd225}: color_data = 12'h800;
			{9'd158, 8'd226}: color_data = 12'h200;
			{9'd158, 8'd227}: color_data = 12'h600;
			{9'd158, 8'd228}: color_data = 12'ha00;
			{9'd158, 8'd229}: color_data = 12'h900;
			{9'd158, 8'd230}: color_data = 12'h300;
			{9'd158, 8'd231}: color_data = 12'h820;
			{9'd158, 8'd232}: color_data = 12'hf30;
			{9'd158, 8'd233}: color_data = 12'hc00;
			{9'd158, 8'd234}: color_data = 12'h500;
			{9'd158, 8'd235}: color_data = 12'h200;
			{9'd158, 8'd236}: color_data = 12'h900;
			{9'd158, 8'd237}: color_data = 12'ha00;
			{9'd158, 8'd238}: color_data = 12'h700;
			{9'd158, 8'd239}: color_data = 12'h100;
			{9'd159, 8'd119}: color_data = 12'h000;
			{9'd159, 8'd120}: color_data = 12'h016;
			{9'd159, 8'd121}: color_data = 12'h017;
			{9'd159, 8'd122}: color_data = 12'h017;
			{9'd159, 8'd123}: color_data = 12'h027;
			{9'd159, 8'd124}: color_data = 12'h027;
			{9'd159, 8'd125}: color_data = 12'h027;
			{9'd159, 8'd126}: color_data = 12'h027;
			{9'd159, 8'd127}: color_data = 12'h028;
			{9'd159, 8'd128}: color_data = 12'h014;
			{9'd159, 8'd129}: color_data = 12'h000;
			{9'd159, 8'd222}: color_data = 12'h300;
			{9'd159, 8'd223}: color_data = 12'hc30;
			{9'd159, 8'd224}: color_data = 12'hc30;
			{9'd159, 8'd225}: color_data = 12'h700;
			{9'd159, 8'd226}: color_data = 12'h100;
			{9'd159, 8'd227}: color_data = 12'h600;
			{9'd159, 8'd228}: color_data = 12'ha00;
			{9'd159, 8'd229}: color_data = 12'h900;
			{9'd159, 8'd230}: color_data = 12'h300;
			{9'd159, 8'd231}: color_data = 12'h620;
			{9'd159, 8'd232}: color_data = 12'hd40;
			{9'd159, 8'd233}: color_data = 12'ha20;
			{9'd159, 8'd234}: color_data = 12'h300;
			{9'd159, 8'd235}: color_data = 12'h200;
			{9'd159, 8'd236}: color_data = 12'h900;
			{9'd159, 8'd237}: color_data = 12'ha00;
			{9'd159, 8'd238}: color_data = 12'h700;
			{9'd159, 8'd239}: color_data = 12'h100;
			{9'd160, 8'd119}: color_data = 12'h000;
			{9'd160, 8'd120}: color_data = 12'h07b;
			{9'd160, 8'd121}: color_data = 12'h0ae;
			{9'd160, 8'd122}: color_data = 12'h09e;
			{9'd160, 8'd123}: color_data = 12'h09e;
			{9'd160, 8'd124}: color_data = 12'h09e;
			{9'd160, 8'd125}: color_data = 12'h09e;
			{9'd160, 8'd126}: color_data = 12'h09e;
			{9'd160, 8'd127}: color_data = 12'h09e;
			{9'd160, 8'd128}: color_data = 12'h057;
			{9'd160, 8'd129}: color_data = 12'h000;
			{9'd160, 8'd222}: color_data = 12'h000;
			{9'd160, 8'd223}: color_data = 12'h200;
			{9'd160, 8'd224}: color_data = 12'h300;
			{9'd160, 8'd225}: color_data = 12'h100;
			{9'd160, 8'd226}: color_data = 12'h000;
			{9'd160, 8'd227}: color_data = 12'h700;
			{9'd160, 8'd228}: color_data = 12'ha00;
			{9'd160, 8'd229}: color_data = 12'h900;
			{9'd160, 8'd230}: color_data = 12'h300;
			{9'd160, 8'd231}: color_data = 12'h100;
			{9'd160, 8'd232}: color_data = 12'h310;
			{9'd160, 8'd233}: color_data = 12'h200;
			{9'd160, 8'd234}: color_data = 12'h000;
			{9'd160, 8'd235}: color_data = 12'h300;
			{9'd160, 8'd236}: color_data = 12'h900;
			{9'd160, 8'd237}: color_data = 12'ha00;
			{9'd160, 8'd238}: color_data = 12'h700;
			{9'd160, 8'd239}: color_data = 12'h100;
			{9'd161, 8'd119}: color_data = 12'h000;
			{9'd161, 8'd120}: color_data = 12'h1ad;
			{9'd161, 8'd121}: color_data = 12'h8ff;
			{9'd161, 8'd122}: color_data = 12'h3df;
			{9'd161, 8'd123}: color_data = 12'h0bf;
			{9'd161, 8'd124}: color_data = 12'h0cf;
			{9'd161, 8'd125}: color_data = 12'h0cf;
			{9'd161, 8'd126}: color_data = 12'h07a;
			{9'd161, 8'd127}: color_data = 12'h08b;
			{9'd161, 8'd128}: color_data = 12'h079;
			{9'd161, 8'd129}: color_data = 12'h000;
			{9'd161, 8'd222}: color_data = 12'h100;
			{9'd161, 8'd223}: color_data = 12'h400;
			{9'd161, 8'd224}: color_data = 12'h500;
			{9'd161, 8'd225}: color_data = 12'h400;
			{9'd161, 8'd226}: color_data = 12'h100;
			{9'd161, 8'd227}: color_data = 12'ha20;
			{9'd161, 8'd228}: color_data = 12'hb10;
			{9'd161, 8'd229}: color_data = 12'h900;
			{9'd161, 8'd230}: color_data = 12'h300;
			{9'd161, 8'd231}: color_data = 12'h200;
			{9'd161, 8'd232}: color_data = 12'h500;
			{9'd161, 8'd233}: color_data = 12'h500;
			{9'd161, 8'd234}: color_data = 12'h200;
			{9'd161, 8'd235}: color_data = 12'h410;
			{9'd161, 8'd236}: color_data = 12'hc20;
			{9'd161, 8'd237}: color_data = 12'ha00;
			{9'd161, 8'd238}: color_data = 12'h700;
			{9'd161, 8'd239}: color_data = 12'h100;
			{9'd162, 8'd119}: color_data = 12'h000;
			{9'd162, 8'd120}: color_data = 12'h2ac;
			{9'd162, 8'd121}: color_data = 12'hdff;
			{9'd162, 8'd122}: color_data = 12'haef;
			{9'd162, 8'd123}: color_data = 12'h1bf;
			{9'd162, 8'd124}: color_data = 12'h0cf;
			{9'd162, 8'd125}: color_data = 12'h08b;
			{9'd162, 8'd126}: color_data = 12'h012;
			{9'd162, 8'd127}: color_data = 12'h068;
			{9'd162, 8'd128}: color_data = 12'h079;
			{9'd162, 8'd129}: color_data = 12'h000;
			{9'd162, 8'd222}: color_data = 12'h200;
			{9'd162, 8'd223}: color_data = 12'h900;
			{9'd162, 8'd224}: color_data = 12'hb00;
			{9'd162, 8'd225}: color_data = 12'h800;
			{9'd162, 8'd226}: color_data = 12'h200;
			{9'd162, 8'd227}: color_data = 12'hb30;
			{9'd162, 8'd228}: color_data = 12'hc10;
			{9'd162, 8'd229}: color_data = 12'h800;
			{9'd162, 8'd230}: color_data = 12'h300;
			{9'd162, 8'd231}: color_data = 12'h400;
			{9'd162, 8'd232}: color_data = 12'ha00;
			{9'd162, 8'd233}: color_data = 12'ha00;
			{9'd162, 8'd234}: color_data = 12'h500;
			{9'd162, 8'd235}: color_data = 12'h510;
			{9'd162, 8'd236}: color_data = 12'hd30;
			{9'd162, 8'd237}: color_data = 12'ha00;
			{9'd162, 8'd238}: color_data = 12'h700;
			{9'd162, 8'd239}: color_data = 12'h100;
			{9'd163, 8'd119}: color_data = 12'h000;
			{9'd163, 8'd120}: color_data = 12'h1ac;
			{9'd163, 8'd121}: color_data = 12'hdff;
			{9'd163, 8'd122}: color_data = 12'hfff;
			{9'd163, 8'd123}: color_data = 12'h8ef;
			{9'd163, 8'd124}: color_data = 12'h19c;
			{9'd163, 8'd125}: color_data = 12'h023;
			{9'd163, 8'd127}: color_data = 12'h068;
			{9'd163, 8'd128}: color_data = 12'h079;
			{9'd163, 8'd129}: color_data = 12'h000;
			{9'd163, 8'd222}: color_data = 12'h200;
			{9'd163, 8'd223}: color_data = 12'h900;
			{9'd163, 8'd224}: color_data = 12'ha00;
			{9'd163, 8'd225}: color_data = 12'h700;
			{9'd163, 8'd226}: color_data = 12'h200;
			{9'd163, 8'd227}: color_data = 12'hb30;
			{9'd163, 8'd228}: color_data = 12'he20;
			{9'd163, 8'd229}: color_data = 12'ha00;
			{9'd163, 8'd230}: color_data = 12'h300;
			{9'd163, 8'd231}: color_data = 12'h400;
			{9'd163, 8'd232}: color_data = 12'ha00;
			{9'd163, 8'd233}: color_data = 12'ha00;
			{9'd163, 8'd234}: color_data = 12'h400;
			{9'd163, 8'd235}: color_data = 12'h510;
			{9'd163, 8'd236}: color_data = 12'hf40;
			{9'd163, 8'd237}: color_data = 12'hd10;
			{9'd163, 8'd238}: color_data = 12'h800;
			{9'd163, 8'd239}: color_data = 12'h100;
			{9'd164, 8'd119}: color_data = 12'h000;
			{9'd164, 8'd120}: color_data = 12'h1ac;
			{9'd164, 8'd121}: color_data = 12'hcff;
			{9'd164, 8'd122}: color_data = 12'hfff;
			{9'd164, 8'd123}: color_data = 12'hddd;
			{9'd164, 8'd124}: color_data = 12'h345;
			{9'd164, 8'd126}: color_data = 12'h000;
			{9'd164, 8'd127}: color_data = 12'h068;
			{9'd164, 8'd128}: color_data = 12'h079;
			{9'd164, 8'd129}: color_data = 12'h000;
			{9'd164, 8'd222}: color_data = 12'h200;
			{9'd164, 8'd223}: color_data = 12'h800;
			{9'd164, 8'd224}: color_data = 12'ha00;
			{9'd164, 8'd225}: color_data = 12'h800;
			{9'd164, 8'd226}: color_data = 12'h200;
			{9'd164, 8'd227}: color_data = 12'h930;
			{9'd164, 8'd228}: color_data = 12'hd30;
			{9'd164, 8'd229}: color_data = 12'h910;
			{9'd164, 8'd230}: color_data = 12'h200;
			{9'd164, 8'd231}: color_data = 12'h400;
			{9'd164, 8'd232}: color_data = 12'h900;
			{9'd164, 8'd233}: color_data = 12'ha00;
			{9'd164, 8'd234}: color_data = 12'h400;
			{9'd164, 8'd235}: color_data = 12'h310;
			{9'd164, 8'd236}: color_data = 12'hc30;
			{9'd164, 8'd237}: color_data = 12'hc20;
			{9'd164, 8'd238}: color_data = 12'h600;
			{9'd164, 8'd239}: color_data = 12'h000;
			{9'd165, 8'd119}: color_data = 12'h000;
			{9'd165, 8'd120}: color_data = 12'h1ac;
			{9'd165, 8'd121}: color_data = 12'hdff;
			{9'd165, 8'd122}: color_data = 12'hfee;
			{9'd165, 8'd123}: color_data = 12'h666;
			{9'd165, 8'd124}: color_data = 12'h002;
			{9'd165, 8'd125}: color_data = 12'h001;
			{9'd165, 8'd126}: color_data = 12'h000;
			{9'd165, 8'd127}: color_data = 12'h068;
			{9'd165, 8'd128}: color_data = 12'h079;
			{9'd165, 8'd129}: color_data = 12'h000;
			{9'd165, 8'd222}: color_data = 12'h200;
			{9'd165, 8'd223}: color_data = 12'h900;
			{9'd165, 8'd224}: color_data = 12'ha00;
			{9'd165, 8'd225}: color_data = 12'h800;
			{9'd165, 8'd226}: color_data = 12'h100;
			{9'd165, 8'd227}: color_data = 12'h100;
			{9'd165, 8'd228}: color_data = 12'h310;
			{9'd165, 8'd229}: color_data = 12'h200;
			{9'd165, 8'd230}: color_data = 12'h000;
			{9'd165, 8'd231}: color_data = 12'h500;
			{9'd165, 8'd232}: color_data = 12'ha00;
			{9'd165, 8'd233}: color_data = 12'ha00;
			{9'd165, 8'd234}: color_data = 12'h500;
			{9'd165, 8'd235}: color_data = 12'h000;
			{9'd165, 8'd236}: color_data = 12'h200;
			{9'd165, 8'd237}: color_data = 12'h300;
			{9'd165, 8'd238}: color_data = 12'h100;
			{9'd165, 8'd239}: color_data = 12'h000;
			{9'd166, 8'd119}: color_data = 12'h000;
			{9'd166, 8'd120}: color_data = 12'h2ad;
			{9'd166, 8'd121}: color_data = 12'hcff;
			{9'd166, 8'd122}: color_data = 12'h877;
			{9'd166, 8'd123}: color_data = 12'h002;
			{9'd166, 8'd124}: color_data = 12'h004;
			{9'd166, 8'd125}: color_data = 12'h004;
			{9'd166, 8'd126}: color_data = 12'h000;
			{9'd166, 8'd127}: color_data = 12'h068;
			{9'd166, 8'd128}: color_data = 12'h079;
			{9'd166, 8'd129}: color_data = 12'h000;
			{9'd166, 8'd222}: color_data = 12'h300;
			{9'd166, 8'd223}: color_data = 12'hc20;
			{9'd166, 8'd224}: color_data = 12'ha00;
			{9'd166, 8'd225}: color_data = 12'h800;
			{9'd166, 8'd226}: color_data = 12'h100;
			{9'd166, 8'd227}: color_data = 12'h300;
			{9'd166, 8'd228}: color_data = 12'h500;
			{9'd166, 8'd229}: color_data = 12'h500;
			{9'd166, 8'd230}: color_data = 12'h100;
			{9'd166, 8'd231}: color_data = 12'h710;
			{9'd166, 8'd232}: color_data = 12'hc10;
			{9'd166, 8'd233}: color_data = 12'h900;
			{9'd166, 8'd234}: color_data = 12'h500;
			{9'd166, 8'd235}: color_data = 12'h100;
			{9'd166, 8'd236}: color_data = 12'h500;
			{9'd166, 8'd237}: color_data = 12'h500;
			{9'd166, 8'd238}: color_data = 12'h400;
			{9'd166, 8'd239}: color_data = 12'h000;
			{9'd167, 8'd119}: color_data = 12'h000;
			{9'd167, 8'd120}: color_data = 12'h1ac;
			{9'd167, 8'd121}: color_data = 12'h689;
			{9'd167, 8'd122}: color_data = 12'h212;
			{9'd167, 8'd123}: color_data = 12'h004;
			{9'd167, 8'd124}: color_data = 12'h005;
			{9'd167, 8'd125}: color_data = 12'h005;
			{9'd167, 8'd126}: color_data = 12'h003;
			{9'd167, 8'd127}: color_data = 12'h06a;
			{9'd167, 8'd128}: color_data = 12'h079;
			{9'd167, 8'd129}: color_data = 12'h000;
			{9'd167, 8'd222}: color_data = 12'h410;
			{9'd167, 8'd223}: color_data = 12'hd30;
			{9'd167, 8'd224}: color_data = 12'hb00;
			{9'd167, 8'd225}: color_data = 12'h700;
			{9'd167, 8'd226}: color_data = 12'h200;
			{9'd167, 8'd227}: color_data = 12'h700;
			{9'd167, 8'd228}: color_data = 12'hb00;
			{9'd167, 8'd229}: color_data = 12'ha00;
			{9'd167, 8'd230}: color_data = 12'h300;
			{9'd167, 8'd231}: color_data = 12'h820;
			{9'd167, 8'd232}: color_data = 12'hd20;
			{9'd167, 8'd233}: color_data = 12'h900;
			{9'd167, 8'd234}: color_data = 12'h500;
			{9'd167, 8'd235}: color_data = 12'h300;
			{9'd167, 8'd236}: color_data = 12'h900;
			{9'd167, 8'd237}: color_data = 12'hb00;
			{9'd167, 8'd238}: color_data = 12'h800;
			{9'd167, 8'd239}: color_data = 12'h100;
			{9'd168, 8'd119}: color_data = 12'h000;
			{9'd168, 8'd120}: color_data = 12'h058;
			{9'd168, 8'd121}: color_data = 12'h013;
			{9'd168, 8'd122}: color_data = 12'h002;
			{9'd168, 8'd123}: color_data = 12'h004;
			{9'd168, 8'd124}: color_data = 12'h004;
			{9'd168, 8'd125}: color_data = 12'h004;
			{9'd168, 8'd126}: color_data = 12'h004;
			{9'd168, 8'd127}: color_data = 12'h038;
			{9'd168, 8'd128}: color_data = 12'h046;
			{9'd168, 8'd129}: color_data = 12'h000;
			{9'd168, 8'd222}: color_data = 12'h410;
			{9'd168, 8'd223}: color_data = 12'he40;
			{9'd168, 8'd224}: color_data = 12'hd20;
			{9'd168, 8'd225}: color_data = 12'h800;
			{9'd168, 8'd226}: color_data = 12'h200;
			{9'd168, 8'd227}: color_data = 12'h600;
			{9'd168, 8'd228}: color_data = 12'ha00;
			{9'd168, 8'd229}: color_data = 12'h900;
			{9'd168, 8'd230}: color_data = 12'h300;
			{9'd168, 8'd231}: color_data = 12'h820;
			{9'd168, 8'd232}: color_data = 12'hf30;
			{9'd168, 8'd233}: color_data = 12'hc00;
			{9'd168, 8'd234}: color_data = 12'h500;
			{9'd168, 8'd235}: color_data = 12'h200;
			{9'd168, 8'd236}: color_data = 12'h900;
			{9'd168, 8'd237}: color_data = 12'ha00;
			{9'd168, 8'd238}: color_data = 12'h700;
			{9'd168, 8'd239}: color_data = 12'h100;
			{9'd169, 8'd119}: color_data = 12'h000;
			{9'd169, 8'd120}: color_data = 12'h016;
			{9'd169, 8'd121}: color_data = 12'h017;
			{9'd169, 8'd122}: color_data = 12'h016;
			{9'd169, 8'd123}: color_data = 12'h027;
			{9'd169, 8'd124}: color_data = 12'h027;
			{9'd169, 8'd125}: color_data = 12'h027;
			{9'd169, 8'd126}: color_data = 12'h027;
			{9'd169, 8'd127}: color_data = 12'h028;
			{9'd169, 8'd128}: color_data = 12'h014;
			{9'd169, 8'd129}: color_data = 12'h000;
			{9'd169, 8'd222}: color_data = 12'h300;
			{9'd169, 8'd223}: color_data = 12'hc30;
			{9'd169, 8'd224}: color_data = 12'hc30;
			{9'd169, 8'd225}: color_data = 12'h700;
			{9'd169, 8'd226}: color_data = 12'h100;
			{9'd169, 8'd227}: color_data = 12'h600;
			{9'd169, 8'd228}: color_data = 12'ha00;
			{9'd169, 8'd229}: color_data = 12'h900;
			{9'd169, 8'd230}: color_data = 12'h300;
			{9'd169, 8'd231}: color_data = 12'h620;
			{9'd169, 8'd232}: color_data = 12'hd40;
			{9'd169, 8'd233}: color_data = 12'ha20;
			{9'd169, 8'd234}: color_data = 12'h300;
			{9'd169, 8'd235}: color_data = 12'h200;
			{9'd169, 8'd236}: color_data = 12'h900;
			{9'd169, 8'd237}: color_data = 12'ha00;
			{9'd169, 8'd238}: color_data = 12'h700;
			{9'd169, 8'd239}: color_data = 12'h100;
			{9'd170, 8'd119}: color_data = 12'h000;
			{9'd170, 8'd120}: color_data = 12'h07b;
			{9'd170, 8'd121}: color_data = 12'h0ae;
			{9'd170, 8'd122}: color_data = 12'h09e;
			{9'd170, 8'd123}: color_data = 12'h09e;
			{9'd170, 8'd124}: color_data = 12'h09e;
			{9'd170, 8'd125}: color_data = 12'h09e;
			{9'd170, 8'd126}: color_data = 12'h09e;
			{9'd170, 8'd127}: color_data = 12'h09e;
			{9'd170, 8'd128}: color_data = 12'h057;
			{9'd170, 8'd129}: color_data = 12'h000;
			{9'd170, 8'd222}: color_data = 12'h000;
			{9'd170, 8'd223}: color_data = 12'h200;
			{9'd170, 8'd224}: color_data = 12'h300;
			{9'd170, 8'd225}: color_data = 12'h100;
			{9'd170, 8'd226}: color_data = 12'h000;
			{9'd170, 8'd227}: color_data = 12'h700;
			{9'd170, 8'd228}: color_data = 12'ha00;
			{9'd170, 8'd229}: color_data = 12'h900;
			{9'd170, 8'd230}: color_data = 12'h300;
			{9'd170, 8'd231}: color_data = 12'h100;
			{9'd170, 8'd232}: color_data = 12'h310;
			{9'd170, 8'd233}: color_data = 12'h200;
			{9'd170, 8'd234}: color_data = 12'h000;
			{9'd170, 8'd235}: color_data = 12'h300;
			{9'd170, 8'd236}: color_data = 12'h900;
			{9'd170, 8'd237}: color_data = 12'ha00;
			{9'd170, 8'd238}: color_data = 12'h700;
			{9'd170, 8'd239}: color_data = 12'h100;
			{9'd171, 8'd119}: color_data = 12'h000;
			{9'd171, 8'd120}: color_data = 12'h1ad;
			{9'd171, 8'd121}: color_data = 12'h8ff;
			{9'd171, 8'd122}: color_data = 12'h3df;
			{9'd171, 8'd123}: color_data = 12'h0cf;
			{9'd171, 8'd124}: color_data = 12'h0cf;
			{9'd171, 8'd125}: color_data = 12'h0cf;
			{9'd171, 8'd126}: color_data = 12'h07a;
			{9'd171, 8'd127}: color_data = 12'h08b;
			{9'd171, 8'd128}: color_data = 12'h079;
			{9'd171, 8'd129}: color_data = 12'h000;
			{9'd171, 8'd222}: color_data = 12'h100;
			{9'd171, 8'd223}: color_data = 12'h500;
			{9'd171, 8'd224}: color_data = 12'h500;
			{9'd171, 8'd225}: color_data = 12'h400;
			{9'd171, 8'd226}: color_data = 12'h200;
			{9'd171, 8'd227}: color_data = 12'ha20;
			{9'd171, 8'd228}: color_data = 12'hb10;
			{9'd171, 8'd229}: color_data = 12'h900;
			{9'd171, 8'd230}: color_data = 12'h300;
			{9'd171, 8'd231}: color_data = 12'h200;
			{9'd171, 8'd232}: color_data = 12'h500;
			{9'd171, 8'd233}: color_data = 12'h500;
			{9'd171, 8'd234}: color_data = 12'h200;
			{9'd171, 8'd235}: color_data = 12'h410;
			{9'd171, 8'd236}: color_data = 12'hc20;
			{9'd171, 8'd237}: color_data = 12'ha00;
			{9'd171, 8'd238}: color_data = 12'h700;
			{9'd171, 8'd239}: color_data = 12'h100;
			{9'd172, 8'd119}: color_data = 12'h000;
			{9'd172, 8'd120}: color_data = 12'h2ac;
			{9'd172, 8'd121}: color_data = 12'hdff;
			{9'd172, 8'd122}: color_data = 12'haef;
			{9'd172, 8'd123}: color_data = 12'h1cf;
			{9'd172, 8'd124}: color_data = 12'h0cf;
			{9'd172, 8'd125}: color_data = 12'h08b;
			{9'd172, 8'd126}: color_data = 12'h012;
			{9'd172, 8'd127}: color_data = 12'h068;
			{9'd172, 8'd128}: color_data = 12'h079;
			{9'd172, 8'd129}: color_data = 12'h000;
			{9'd172, 8'd222}: color_data = 12'h200;
			{9'd172, 8'd223}: color_data = 12'h900;
			{9'd172, 8'd224}: color_data = 12'hb00;
			{9'd172, 8'd225}: color_data = 12'h800;
			{9'd172, 8'd226}: color_data = 12'h200;
			{9'd172, 8'd227}: color_data = 12'hb30;
			{9'd172, 8'd228}: color_data = 12'hc10;
			{9'd172, 8'd229}: color_data = 12'h800;
			{9'd172, 8'd230}: color_data = 12'h300;
			{9'd172, 8'd231}: color_data = 12'h400;
			{9'd172, 8'd232}: color_data = 12'ha00;
			{9'd172, 8'd233}: color_data = 12'ha00;
			{9'd172, 8'd234}: color_data = 12'h500;
			{9'd172, 8'd235}: color_data = 12'h510;
			{9'd172, 8'd236}: color_data = 12'hd30;
			{9'd172, 8'd237}: color_data = 12'ha00;
			{9'd172, 8'd238}: color_data = 12'h700;
			{9'd172, 8'd239}: color_data = 12'h100;
			{9'd173, 8'd119}: color_data = 12'h000;
			{9'd173, 8'd120}: color_data = 12'h1ac;
			{9'd173, 8'd121}: color_data = 12'hdff;
			{9'd173, 8'd122}: color_data = 12'hfff;
			{9'd173, 8'd123}: color_data = 12'h8ef;
			{9'd173, 8'd124}: color_data = 12'h19c;
			{9'd173, 8'd125}: color_data = 12'h023;
			{9'd173, 8'd127}: color_data = 12'h068;
			{9'd173, 8'd128}: color_data = 12'h079;
			{9'd173, 8'd129}: color_data = 12'h000;
			{9'd173, 8'd222}: color_data = 12'h200;
			{9'd173, 8'd223}: color_data = 12'h900;
			{9'd173, 8'd224}: color_data = 12'ha00;
			{9'd173, 8'd225}: color_data = 12'h700;
			{9'd173, 8'd226}: color_data = 12'h200;
			{9'd173, 8'd227}: color_data = 12'hb30;
			{9'd173, 8'd228}: color_data = 12'he20;
			{9'd173, 8'd229}: color_data = 12'ha00;
			{9'd173, 8'd230}: color_data = 12'h300;
			{9'd173, 8'd231}: color_data = 12'h400;
			{9'd173, 8'd232}: color_data = 12'ha00;
			{9'd173, 8'd233}: color_data = 12'ha00;
			{9'd173, 8'd234}: color_data = 12'h400;
			{9'd173, 8'd235}: color_data = 12'h510;
			{9'd173, 8'd236}: color_data = 12'hf40;
			{9'd173, 8'd237}: color_data = 12'hd10;
			{9'd173, 8'd238}: color_data = 12'h800;
			{9'd173, 8'd239}: color_data = 12'h100;
			{9'd174, 8'd119}: color_data = 12'h000;
			{9'd174, 8'd120}: color_data = 12'h1ac;
			{9'd174, 8'd121}: color_data = 12'hcff;
			{9'd174, 8'd122}: color_data = 12'hfff;
			{9'd174, 8'd123}: color_data = 12'hddd;
			{9'd174, 8'd124}: color_data = 12'h345;
			{9'd174, 8'd126}: color_data = 12'h000;
			{9'd174, 8'd127}: color_data = 12'h068;
			{9'd174, 8'd128}: color_data = 12'h079;
			{9'd174, 8'd129}: color_data = 12'h000;
			{9'd174, 8'd222}: color_data = 12'h200;
			{9'd174, 8'd223}: color_data = 12'h800;
			{9'd174, 8'd224}: color_data = 12'ha00;
			{9'd174, 8'd225}: color_data = 12'h800;
			{9'd174, 8'd226}: color_data = 12'h200;
			{9'd174, 8'd227}: color_data = 12'h920;
			{9'd174, 8'd228}: color_data = 12'hd30;
			{9'd174, 8'd229}: color_data = 12'h910;
			{9'd174, 8'd230}: color_data = 12'h200;
			{9'd174, 8'd231}: color_data = 12'h400;
			{9'd174, 8'd232}: color_data = 12'h900;
			{9'd174, 8'd233}: color_data = 12'ha00;
			{9'd174, 8'd234}: color_data = 12'h400;
			{9'd174, 8'd235}: color_data = 12'h310;
			{9'd174, 8'd236}: color_data = 12'hc30;
			{9'd174, 8'd237}: color_data = 12'hc20;
			{9'd174, 8'd238}: color_data = 12'h600;
			{9'd174, 8'd239}: color_data = 12'h000;
			{9'd175, 8'd119}: color_data = 12'h000;
			{9'd175, 8'd120}: color_data = 12'h1ac;
			{9'd175, 8'd121}: color_data = 12'hdff;
			{9'd175, 8'd122}: color_data = 12'hfee;
			{9'd175, 8'd123}: color_data = 12'h666;
			{9'd175, 8'd124}: color_data = 12'h002;
			{9'd175, 8'd125}: color_data = 12'h001;
			{9'd175, 8'd126}: color_data = 12'h000;
			{9'd175, 8'd127}: color_data = 12'h068;
			{9'd175, 8'd128}: color_data = 12'h079;
			{9'd175, 8'd129}: color_data = 12'h000;
			{9'd175, 8'd222}: color_data = 12'h200;
			{9'd175, 8'd223}: color_data = 12'h900;
			{9'd175, 8'd224}: color_data = 12'ha00;
			{9'd175, 8'd225}: color_data = 12'h800;
			{9'd175, 8'd226}: color_data = 12'h100;
			{9'd175, 8'd227}: color_data = 12'h100;
			{9'd175, 8'd228}: color_data = 12'h310;
			{9'd175, 8'd229}: color_data = 12'h200;
			{9'd175, 8'd230}: color_data = 12'h000;
			{9'd175, 8'd231}: color_data = 12'h500;
			{9'd175, 8'd232}: color_data = 12'ha00;
			{9'd175, 8'd233}: color_data = 12'ha00;
			{9'd175, 8'd234}: color_data = 12'h500;
			{9'd175, 8'd235}: color_data = 12'h000;
			{9'd175, 8'd236}: color_data = 12'h200;
			{9'd175, 8'd237}: color_data = 12'h300;
			{9'd175, 8'd238}: color_data = 12'h100;
			{9'd175, 8'd239}: color_data = 12'h000;
			{9'd176, 8'd119}: color_data = 12'h000;
			{9'd176, 8'd120}: color_data = 12'h2ad;
			{9'd176, 8'd121}: color_data = 12'hcff;
			{9'd176, 8'd122}: color_data = 12'h877;
			{9'd176, 8'd123}: color_data = 12'h002;
			{9'd176, 8'd124}: color_data = 12'h004;
			{9'd176, 8'd125}: color_data = 12'h004;
			{9'd176, 8'd126}: color_data = 12'h000;
			{9'd176, 8'd127}: color_data = 12'h068;
			{9'd176, 8'd128}: color_data = 12'h079;
			{9'd176, 8'd129}: color_data = 12'h000;
			{9'd176, 8'd222}: color_data = 12'h300;
			{9'd176, 8'd223}: color_data = 12'hc20;
			{9'd176, 8'd224}: color_data = 12'ha00;
			{9'd176, 8'd225}: color_data = 12'h800;
			{9'd176, 8'd226}: color_data = 12'h100;
			{9'd176, 8'd227}: color_data = 12'h300;
			{9'd176, 8'd228}: color_data = 12'h500;
			{9'd176, 8'd229}: color_data = 12'h500;
			{9'd176, 8'd230}: color_data = 12'h100;
			{9'd176, 8'd231}: color_data = 12'h710;
			{9'd176, 8'd232}: color_data = 12'hc10;
			{9'd176, 8'd233}: color_data = 12'h900;
			{9'd176, 8'd234}: color_data = 12'h500;
			{9'd176, 8'd235}: color_data = 12'h100;
			{9'd176, 8'd236}: color_data = 12'h500;
			{9'd176, 8'd237}: color_data = 12'h600;
			{9'd176, 8'd238}: color_data = 12'h400;
			{9'd176, 8'd239}: color_data = 12'h000;
			{9'd177, 8'd119}: color_data = 12'h000;
			{9'd177, 8'd120}: color_data = 12'h1ac;
			{9'd177, 8'd121}: color_data = 12'h689;
			{9'd177, 8'd122}: color_data = 12'h212;
			{9'd177, 8'd123}: color_data = 12'h004;
			{9'd177, 8'd124}: color_data = 12'h005;
			{9'd177, 8'd125}: color_data = 12'h005;
			{9'd177, 8'd126}: color_data = 12'h003;
			{9'd177, 8'd127}: color_data = 12'h06a;
			{9'd177, 8'd128}: color_data = 12'h079;
			{9'd177, 8'd129}: color_data = 12'h000;
			{9'd177, 8'd222}: color_data = 12'h410;
			{9'd177, 8'd223}: color_data = 12'hd30;
			{9'd177, 8'd224}: color_data = 12'hb00;
			{9'd177, 8'd225}: color_data = 12'h700;
			{9'd177, 8'd226}: color_data = 12'h200;
			{9'd177, 8'd227}: color_data = 12'h700;
			{9'd177, 8'd228}: color_data = 12'hb00;
			{9'd177, 8'd229}: color_data = 12'h900;
			{9'd177, 8'd230}: color_data = 12'h300;
			{9'd177, 8'd231}: color_data = 12'h820;
			{9'd177, 8'd232}: color_data = 12'hd20;
			{9'd177, 8'd233}: color_data = 12'h900;
			{9'd177, 8'd234}: color_data = 12'h500;
			{9'd177, 8'd235}: color_data = 12'h300;
			{9'd177, 8'd236}: color_data = 12'h900;
			{9'd177, 8'd237}: color_data = 12'hb00;
			{9'd177, 8'd238}: color_data = 12'h800;
			{9'd177, 8'd239}: color_data = 12'h100;
			{9'd178, 8'd119}: color_data = 12'h000;
			{9'd178, 8'd120}: color_data = 12'h058;
			{9'd178, 8'd121}: color_data = 12'h013;
			{9'd178, 8'd122}: color_data = 12'h002;
			{9'd178, 8'd123}: color_data = 12'h004;
			{9'd178, 8'd124}: color_data = 12'h004;
			{9'd178, 8'd125}: color_data = 12'h004;
			{9'd178, 8'd126}: color_data = 12'h004;
			{9'd178, 8'd127}: color_data = 12'h038;
			{9'd178, 8'd128}: color_data = 12'h046;
			{9'd178, 8'd129}: color_data = 12'h000;
			{9'd178, 8'd222}: color_data = 12'h410;
			{9'd178, 8'd223}: color_data = 12'he40;
			{9'd178, 8'd224}: color_data = 12'hd20;
			{9'd178, 8'd225}: color_data = 12'h800;
			{9'd178, 8'd226}: color_data = 12'h200;
			{9'd178, 8'd227}: color_data = 12'h600;
			{9'd178, 8'd228}: color_data = 12'ha00;
			{9'd178, 8'd229}: color_data = 12'h900;
			{9'd178, 8'd230}: color_data = 12'h300;
			{9'd178, 8'd231}: color_data = 12'h820;
			{9'd178, 8'd232}: color_data = 12'hf30;
			{9'd178, 8'd233}: color_data = 12'hc00;
			{9'd178, 8'd234}: color_data = 12'h500;
			{9'd178, 8'd235}: color_data = 12'h200;
			{9'd178, 8'd236}: color_data = 12'h900;
			{9'd178, 8'd237}: color_data = 12'ha00;
			{9'd178, 8'd238}: color_data = 12'h700;
			{9'd178, 8'd239}: color_data = 12'h100;
			{9'd179, 8'd68}: color_data = 12'h001;
			{9'd179, 8'd69}: color_data = 12'h023;
			{9'd179, 8'd70}: color_data = 12'h012;
			{9'd179, 8'd71}: color_data = 12'h022;
			{9'd179, 8'd72}: color_data = 12'h022;
			{9'd179, 8'd73}: color_data = 12'h022;
			{9'd179, 8'd74}: color_data = 12'h023;
			{9'd179, 8'd75}: color_data = 12'h023;
			{9'd179, 8'd76}: color_data = 12'h022;
			{9'd179, 8'd77}: color_data = 12'h000;
			{9'd179, 8'd119}: color_data = 12'h000;
			{9'd179, 8'd120}: color_data = 12'h016;
			{9'd179, 8'd121}: color_data = 12'h027;
			{9'd179, 8'd122}: color_data = 12'h026;
			{9'd179, 8'd123}: color_data = 12'h027;
			{9'd179, 8'd124}: color_data = 12'h027;
			{9'd179, 8'd125}: color_data = 12'h027;
			{9'd179, 8'd126}: color_data = 12'h027;
			{9'd179, 8'd127}: color_data = 12'h028;
			{9'd179, 8'd128}: color_data = 12'h014;
			{9'd179, 8'd129}: color_data = 12'h000;
			{9'd179, 8'd222}: color_data = 12'h300;
			{9'd179, 8'd223}: color_data = 12'hc30;
			{9'd179, 8'd224}: color_data = 12'hc30;
			{9'd179, 8'd225}: color_data = 12'h600;
			{9'd179, 8'd226}: color_data = 12'h100;
			{9'd179, 8'd227}: color_data = 12'h600;
			{9'd179, 8'd228}: color_data = 12'ha00;
			{9'd179, 8'd229}: color_data = 12'h900;
			{9'd179, 8'd230}: color_data = 12'h300;
			{9'd179, 8'd231}: color_data = 12'h620;
			{9'd179, 8'd232}: color_data = 12'hd40;
			{9'd179, 8'd233}: color_data = 12'ha20;
			{9'd179, 8'd234}: color_data = 12'h300;
			{9'd179, 8'd235}: color_data = 12'h200;
			{9'd179, 8'd236}: color_data = 12'h900;
			{9'd179, 8'd237}: color_data = 12'ha00;
			{9'd179, 8'd238}: color_data = 12'h700;
			{9'd179, 8'd239}: color_data = 12'h100;
			{9'd180, 8'd68}: color_data = 12'h045;
			{9'd180, 8'd69}: color_data = 12'h0ad;
			{9'd180, 8'd70}: color_data = 12'h09d;
			{9'd180, 8'd71}: color_data = 12'h09d;
			{9'd180, 8'd72}: color_data = 12'h09d;
			{9'd180, 8'd73}: color_data = 12'h09d;
			{9'd180, 8'd74}: color_data = 12'h09d;
			{9'd180, 8'd75}: color_data = 12'h09d;
			{9'd180, 8'd76}: color_data = 12'h09c;
			{9'd180, 8'd77}: color_data = 12'h023;
			{9'd180, 8'd119}: color_data = 12'h000;
			{9'd180, 8'd120}: color_data = 12'h07b;
			{9'd180, 8'd121}: color_data = 12'h0ae;
			{9'd180, 8'd122}: color_data = 12'h09e;
			{9'd180, 8'd123}: color_data = 12'h09e;
			{9'd180, 8'd124}: color_data = 12'h09e;
			{9'd180, 8'd125}: color_data = 12'h09e;
			{9'd180, 8'd126}: color_data = 12'h09e;
			{9'd180, 8'd127}: color_data = 12'h09e;
			{9'd180, 8'd128}: color_data = 12'h057;
			{9'd180, 8'd129}: color_data = 12'h000;
			{9'd180, 8'd222}: color_data = 12'h000;
			{9'd180, 8'd223}: color_data = 12'h200;
			{9'd180, 8'd224}: color_data = 12'h300;
			{9'd180, 8'd225}: color_data = 12'h100;
			{9'd180, 8'd226}: color_data = 12'h000;
			{9'd180, 8'd227}: color_data = 12'h700;
			{9'd180, 8'd228}: color_data = 12'ha00;
			{9'd180, 8'd229}: color_data = 12'h900;
			{9'd180, 8'd230}: color_data = 12'h300;
			{9'd180, 8'd231}: color_data = 12'h100;
			{9'd180, 8'd232}: color_data = 12'h310;
			{9'd180, 8'd233}: color_data = 12'h200;
			{9'd180, 8'd234}: color_data = 12'h000;
			{9'd180, 8'd235}: color_data = 12'h300;
			{9'd180, 8'd236}: color_data = 12'h900;
			{9'd180, 8'd237}: color_data = 12'ha00;
			{9'd180, 8'd238}: color_data = 12'h700;
			{9'd180, 8'd239}: color_data = 12'h100;
			{9'd181, 8'd68}: color_data = 12'h057;
			{9'd181, 8'd69}: color_data = 12'h4ef;
			{9'd181, 8'd70}: color_data = 12'h7ef;
			{9'd181, 8'd71}: color_data = 12'h0cf;
			{9'd181, 8'd72}: color_data = 12'h0cf;
			{9'd181, 8'd73}: color_data = 12'h0df;
			{9'd181, 8'd74}: color_data = 12'h0be;
			{9'd181, 8'd75}: color_data = 12'h069;
			{9'd181, 8'd76}: color_data = 12'h09d;
			{9'd181, 8'd77}: color_data = 12'h034;
			{9'd181, 8'd119}: color_data = 12'h000;
			{9'd181, 8'd120}: color_data = 12'h1ad;
			{9'd181, 8'd121}: color_data = 12'h8ff;
			{9'd181, 8'd122}: color_data = 12'h3df;
			{9'd181, 8'd123}: color_data = 12'h0bf;
			{9'd181, 8'd124}: color_data = 12'h0cf;
			{9'd181, 8'd125}: color_data = 12'h0cf;
			{9'd181, 8'd126}: color_data = 12'h079;
			{9'd181, 8'd127}: color_data = 12'h08b;
			{9'd181, 8'd128}: color_data = 12'h079;
			{9'd181, 8'd129}: color_data = 12'h000;
			{9'd181, 8'd222}: color_data = 12'h100;
			{9'd181, 8'd223}: color_data = 12'h500;
			{9'd181, 8'd224}: color_data = 12'h500;
			{9'd181, 8'd225}: color_data = 12'h400;
			{9'd181, 8'd226}: color_data = 12'h100;
			{9'd181, 8'd227}: color_data = 12'ha20;
			{9'd181, 8'd228}: color_data = 12'hb10;
			{9'd181, 8'd229}: color_data = 12'h900;
			{9'd181, 8'd230}: color_data = 12'h300;
			{9'd181, 8'd231}: color_data = 12'h200;
			{9'd181, 8'd232}: color_data = 12'h500;
			{9'd181, 8'd233}: color_data = 12'h500;
			{9'd181, 8'd234}: color_data = 12'h200;
			{9'd181, 8'd235}: color_data = 12'h410;
			{9'd181, 8'd236}: color_data = 12'hc20;
			{9'd181, 8'd237}: color_data = 12'ha00;
			{9'd181, 8'd238}: color_data = 12'h700;
			{9'd181, 8'd239}: color_data = 12'h100;
			{9'd182, 8'd68}: color_data = 12'h047;
			{9'd182, 8'd69}: color_data = 12'h6df;
			{9'd182, 8'd70}: color_data = 12'heff;
			{9'd182, 8'd71}: color_data = 12'h6df;
			{9'd182, 8'd72}: color_data = 12'h0bf;
			{9'd182, 8'd73}: color_data = 12'h0bf;
			{9'd182, 8'd74}: color_data = 12'h056;
			{9'd182, 8'd75}: color_data = 12'h012;
			{9'd182, 8'd76}: color_data = 12'h08b;
			{9'd182, 8'd77}: color_data = 12'h034;
			{9'd182, 8'd119}: color_data = 12'h000;
			{9'd182, 8'd120}: color_data = 12'h2ac;
			{9'd182, 8'd121}: color_data = 12'hdff;
			{9'd182, 8'd122}: color_data = 12'haef;
			{9'd182, 8'd123}: color_data = 12'h1cf;
			{9'd182, 8'd124}: color_data = 12'h0cf;
			{9'd182, 8'd125}: color_data = 12'h08b;
			{9'd182, 8'd126}: color_data = 12'h012;
			{9'd182, 8'd127}: color_data = 12'h068;
			{9'd182, 8'd128}: color_data = 12'h079;
			{9'd182, 8'd129}: color_data = 12'h000;
			{9'd182, 8'd222}: color_data = 12'h200;
			{9'd182, 8'd223}: color_data = 12'h900;
			{9'd182, 8'd224}: color_data = 12'hb00;
			{9'd182, 8'd225}: color_data = 12'h800;
			{9'd182, 8'd226}: color_data = 12'h200;
			{9'd182, 8'd227}: color_data = 12'hb30;
			{9'd182, 8'd228}: color_data = 12'hc10;
			{9'd182, 8'd229}: color_data = 12'h800;
			{9'd182, 8'd230}: color_data = 12'h300;
			{9'd182, 8'd231}: color_data = 12'h500;
			{9'd182, 8'd232}: color_data = 12'ha00;
			{9'd182, 8'd233}: color_data = 12'ha00;
			{9'd182, 8'd234}: color_data = 12'h500;
			{9'd182, 8'd235}: color_data = 12'h510;
			{9'd182, 8'd236}: color_data = 12'hd30;
			{9'd182, 8'd237}: color_data = 12'ha00;
			{9'd182, 8'd238}: color_data = 12'h700;
			{9'd182, 8'd239}: color_data = 12'h100;
			{9'd183, 8'd68}: color_data = 12'h047;
			{9'd183, 8'd69}: color_data = 12'h6df;
			{9'd183, 8'd70}: color_data = 12'hfff;
			{9'd183, 8'd71}: color_data = 12'hdff;
			{9'd183, 8'd72}: color_data = 12'h5df;
			{9'd183, 8'd73}: color_data = 12'h068;
			{9'd183, 8'd74}: color_data = 12'h000;
			{9'd183, 8'd75}: color_data = 12'h012;
			{9'd183, 8'd76}: color_data = 12'h08c;
			{9'd183, 8'd77}: color_data = 12'h034;
			{9'd183, 8'd119}: color_data = 12'h000;
			{9'd183, 8'd120}: color_data = 12'h1ac;
			{9'd183, 8'd121}: color_data = 12'hdff;
			{9'd183, 8'd122}: color_data = 12'hfff;
			{9'd183, 8'd123}: color_data = 12'h8ef;
			{9'd183, 8'd124}: color_data = 12'h19c;
			{9'd183, 8'd125}: color_data = 12'h023;
			{9'd183, 8'd127}: color_data = 12'h068;
			{9'd183, 8'd128}: color_data = 12'h079;
			{9'd183, 8'd129}: color_data = 12'h000;
			{9'd183, 8'd222}: color_data = 12'h200;
			{9'd183, 8'd223}: color_data = 12'h900;
			{9'd183, 8'd224}: color_data = 12'ha00;
			{9'd183, 8'd225}: color_data = 12'h700;
			{9'd183, 8'd226}: color_data = 12'h200;
			{9'd183, 8'd227}: color_data = 12'hb30;
			{9'd183, 8'd228}: color_data = 12'he20;
			{9'd183, 8'd229}: color_data = 12'ha00;
			{9'd183, 8'd230}: color_data = 12'h300;
			{9'd183, 8'd231}: color_data = 12'h400;
			{9'd183, 8'd232}: color_data = 12'ha00;
			{9'd183, 8'd233}: color_data = 12'ha00;
			{9'd183, 8'd234}: color_data = 12'h400;
			{9'd183, 8'd235}: color_data = 12'h510;
			{9'd183, 8'd236}: color_data = 12'hf40;
			{9'd183, 8'd237}: color_data = 12'hd10;
			{9'd183, 8'd238}: color_data = 12'h800;
			{9'd183, 8'd239}: color_data = 12'h100;
			{9'd184, 8'd68}: color_data = 12'h047;
			{9'd184, 8'd69}: color_data = 12'h6df;
			{9'd184, 8'd70}: color_data = 12'hfff;
			{9'd184, 8'd71}: color_data = 12'hfff;
			{9'd184, 8'd72}: color_data = 12'h9aa;
			{9'd184, 8'd73}: color_data = 12'h011;
			{9'd184, 8'd75}: color_data = 12'h012;
			{9'd184, 8'd76}: color_data = 12'h08c;
			{9'd184, 8'd77}: color_data = 12'h034;
			{9'd184, 8'd119}: color_data = 12'h000;
			{9'd184, 8'd120}: color_data = 12'h1ac;
			{9'd184, 8'd121}: color_data = 12'hcff;
			{9'd184, 8'd122}: color_data = 12'hfff;
			{9'd184, 8'd123}: color_data = 12'hddd;
			{9'd184, 8'd124}: color_data = 12'h345;
			{9'd184, 8'd126}: color_data = 12'h000;
			{9'd184, 8'd127}: color_data = 12'h068;
			{9'd184, 8'd128}: color_data = 12'h079;
			{9'd184, 8'd129}: color_data = 12'h000;
			{9'd184, 8'd222}: color_data = 12'h200;
			{9'd184, 8'd223}: color_data = 12'h800;
			{9'd184, 8'd224}: color_data = 12'ha00;
			{9'd184, 8'd225}: color_data = 12'h700;
			{9'd184, 8'd226}: color_data = 12'h200;
			{9'd184, 8'd227}: color_data = 12'h920;
			{9'd184, 8'd228}: color_data = 12'hd30;
			{9'd184, 8'd229}: color_data = 12'h910;
			{9'd184, 8'd230}: color_data = 12'h200;
			{9'd184, 8'd231}: color_data = 12'h400;
			{9'd184, 8'd232}: color_data = 12'h900;
			{9'd184, 8'd233}: color_data = 12'ha00;
			{9'd184, 8'd234}: color_data = 12'h400;
			{9'd184, 8'd235}: color_data = 12'h310;
			{9'd184, 8'd236}: color_data = 12'hc30;
			{9'd184, 8'd237}: color_data = 12'hc20;
			{9'd184, 8'd238}: color_data = 12'h600;
			{9'd184, 8'd239}: color_data = 12'h000;
			{9'd185, 8'd68}: color_data = 12'h047;
			{9'd185, 8'd69}: color_data = 12'h6df;
			{9'd185, 8'd70}: color_data = 12'hfff;
			{9'd185, 8'd71}: color_data = 12'hcbb;
			{9'd185, 8'd72}: color_data = 12'h323;
			{9'd185, 8'd73}: color_data = 12'h002;
			{9'd185, 8'd74}: color_data = 12'h000;
			{9'd185, 8'd75}: color_data = 12'h012;
			{9'd185, 8'd76}: color_data = 12'h08c;
			{9'd185, 8'd77}: color_data = 12'h034;
			{9'd185, 8'd119}: color_data = 12'h000;
			{9'd185, 8'd120}: color_data = 12'h1ac;
			{9'd185, 8'd121}: color_data = 12'hdff;
			{9'd185, 8'd122}: color_data = 12'hfee;
			{9'd185, 8'd123}: color_data = 12'h666;
			{9'd185, 8'd124}: color_data = 12'h002;
			{9'd185, 8'd125}: color_data = 12'h001;
			{9'd185, 8'd126}: color_data = 12'h000;
			{9'd185, 8'd127}: color_data = 12'h068;
			{9'd185, 8'd128}: color_data = 12'h079;
			{9'd185, 8'd129}: color_data = 12'h000;
			{9'd185, 8'd222}: color_data = 12'h200;
			{9'd185, 8'd223}: color_data = 12'h900;
			{9'd185, 8'd224}: color_data = 12'ha00;
			{9'd185, 8'd225}: color_data = 12'h800;
			{9'd185, 8'd226}: color_data = 12'h100;
			{9'd185, 8'd227}: color_data = 12'h100;
			{9'd185, 8'd228}: color_data = 12'h310;
			{9'd185, 8'd229}: color_data = 12'h200;
			{9'd185, 8'd230}: color_data = 12'h000;
			{9'd185, 8'd231}: color_data = 12'h500;
			{9'd185, 8'd232}: color_data = 12'ha00;
			{9'd185, 8'd233}: color_data = 12'ha00;
			{9'd185, 8'd234}: color_data = 12'h500;
			{9'd185, 8'd235}: color_data = 12'h000;
			{9'd185, 8'd236}: color_data = 12'h200;
			{9'd185, 8'd237}: color_data = 12'h300;
			{9'd185, 8'd238}: color_data = 12'h100;
			{9'd185, 8'd239}: color_data = 12'h000;
			{9'd186, 8'd68}: color_data = 12'h047;
			{9'd186, 8'd69}: color_data = 12'h6ef;
			{9'd186, 8'd70}: color_data = 12'hddc;
			{9'd186, 8'd71}: color_data = 12'h434;
			{9'd186, 8'd72}: color_data = 12'h003;
			{9'd186, 8'd73}: color_data = 12'h005;
			{9'd186, 8'd74}: color_data = 12'h002;
			{9'd186, 8'd75}: color_data = 12'h012;
			{9'd186, 8'd76}: color_data = 12'h08c;
			{9'd186, 8'd77}: color_data = 12'h034;
			{9'd186, 8'd119}: color_data = 12'h000;
			{9'd186, 8'd120}: color_data = 12'h2ad;
			{9'd186, 8'd121}: color_data = 12'hcff;
			{9'd186, 8'd122}: color_data = 12'h877;
			{9'd186, 8'd123}: color_data = 12'h002;
			{9'd186, 8'd124}: color_data = 12'h004;
			{9'd186, 8'd125}: color_data = 12'h004;
			{9'd186, 8'd126}: color_data = 12'h000;
			{9'd186, 8'd127}: color_data = 12'h068;
			{9'd186, 8'd128}: color_data = 12'h079;
			{9'd186, 8'd129}: color_data = 12'h000;
			{9'd186, 8'd222}: color_data = 12'h300;
			{9'd186, 8'd223}: color_data = 12'hc20;
			{9'd186, 8'd224}: color_data = 12'ha00;
			{9'd186, 8'd225}: color_data = 12'h800;
			{9'd186, 8'd226}: color_data = 12'h200;
			{9'd186, 8'd227}: color_data = 12'h300;
			{9'd186, 8'd228}: color_data = 12'h500;
			{9'd186, 8'd229}: color_data = 12'h500;
			{9'd186, 8'd230}: color_data = 12'h100;
			{9'd186, 8'd231}: color_data = 12'h710;
			{9'd186, 8'd232}: color_data = 12'hc10;
			{9'd186, 8'd233}: color_data = 12'h900;
			{9'd186, 8'd234}: color_data = 12'h500;
			{9'd186, 8'd235}: color_data = 12'h100;
			{9'd186, 8'd236}: color_data = 12'h500;
			{9'd186, 8'd237}: color_data = 12'h500;
			{9'd186, 8'd238}: color_data = 12'h400;
			{9'd186, 8'd239}: color_data = 12'h000;
			{9'd187, 8'd68}: color_data = 12'h057;
			{9'd187, 8'd69}: color_data = 12'h3bd;
			{9'd187, 8'd70}: color_data = 12'h555;
			{9'd187, 8'd71}: color_data = 12'h002;
			{9'd187, 8'd72}: color_data = 12'h005;
			{9'd187, 8'd73}: color_data = 12'h005;
			{9'd187, 8'd74}: color_data = 12'h004;
			{9'd187, 8'd75}: color_data = 12'h025;
			{9'd187, 8'd76}: color_data = 12'h09c;
			{9'd187, 8'd77}: color_data = 12'h034;
			{9'd187, 8'd119}: color_data = 12'h000;
			{9'd187, 8'd120}: color_data = 12'h1ac;
			{9'd187, 8'd121}: color_data = 12'h689;
			{9'd187, 8'd122}: color_data = 12'h212;
			{9'd187, 8'd123}: color_data = 12'h004;
			{9'd187, 8'd124}: color_data = 12'h005;
			{9'd187, 8'd125}: color_data = 12'h005;
			{9'd187, 8'd126}: color_data = 12'h003;
			{9'd187, 8'd127}: color_data = 12'h06a;
			{9'd187, 8'd128}: color_data = 12'h079;
			{9'd187, 8'd129}: color_data = 12'h000;
			{9'd187, 8'd222}: color_data = 12'h410;
			{9'd187, 8'd223}: color_data = 12'hd30;
			{9'd187, 8'd224}: color_data = 12'hb00;
			{9'd187, 8'd225}: color_data = 12'h700;
			{9'd187, 8'd226}: color_data = 12'h200;
			{9'd187, 8'd227}: color_data = 12'h700;
			{9'd187, 8'd228}: color_data = 12'hb00;
			{9'd187, 8'd229}: color_data = 12'ha00;
			{9'd187, 8'd230}: color_data = 12'h300;
			{9'd187, 8'd231}: color_data = 12'h820;
			{9'd187, 8'd232}: color_data = 12'hd20;
			{9'd187, 8'd233}: color_data = 12'h900;
			{9'd187, 8'd234}: color_data = 12'h500;
			{9'd187, 8'd235}: color_data = 12'h300;
			{9'd187, 8'd236}: color_data = 12'h900;
			{9'd187, 8'd237}: color_data = 12'hb00;
			{9'd187, 8'd238}: color_data = 12'h800;
			{9'd187, 8'd239}: color_data = 12'h100;
			{9'd188, 8'd68}: color_data = 12'h035;
			{9'd188, 8'd69}: color_data = 12'h047;
			{9'd188, 8'd70}: color_data = 12'h001;
			{9'd188, 8'd71}: color_data = 12'h004;
			{9'd188, 8'd72}: color_data = 12'h004;
			{9'd188, 8'd73}: color_data = 12'h004;
			{9'd188, 8'd74}: color_data = 12'h004;
			{9'd188, 8'd75}: color_data = 12'h015;
			{9'd188, 8'd76}: color_data = 12'h059;
			{9'd188, 8'd77}: color_data = 12'h023;
			{9'd188, 8'd119}: color_data = 12'h000;
			{9'd188, 8'd120}: color_data = 12'h058;
			{9'd188, 8'd121}: color_data = 12'h013;
			{9'd188, 8'd122}: color_data = 12'h002;
			{9'd188, 8'd123}: color_data = 12'h004;
			{9'd188, 8'd124}: color_data = 12'h004;
			{9'd188, 8'd125}: color_data = 12'h004;
			{9'd188, 8'd126}: color_data = 12'h004;
			{9'd188, 8'd127}: color_data = 12'h039;
			{9'd188, 8'd128}: color_data = 12'h046;
			{9'd188, 8'd129}: color_data = 12'h000;
			{9'd188, 8'd222}: color_data = 12'h410;
			{9'd188, 8'd223}: color_data = 12'he40;
			{9'd188, 8'd224}: color_data = 12'hd20;
			{9'd188, 8'd225}: color_data = 12'h800;
			{9'd188, 8'd226}: color_data = 12'h200;
			{9'd188, 8'd227}: color_data = 12'h600;
			{9'd188, 8'd228}: color_data = 12'ha00;
			{9'd188, 8'd229}: color_data = 12'h900;
			{9'd188, 8'd230}: color_data = 12'h300;
			{9'd188, 8'd231}: color_data = 12'h820;
			{9'd188, 8'd232}: color_data = 12'hf30;
			{9'd188, 8'd233}: color_data = 12'hc00;
			{9'd188, 8'd234}: color_data = 12'h500;
			{9'd188, 8'd235}: color_data = 12'h200;
			{9'd188, 8'd236}: color_data = 12'h900;
			{9'd188, 8'd237}: color_data = 12'ha00;
			{9'd188, 8'd238}: color_data = 12'h700;
			{9'd188, 8'd239}: color_data = 12'h100;
			{9'd189, 8'd68}: color_data = 12'h013;
			{9'd189, 8'd69}: color_data = 12'h027;
			{9'd189, 8'd70}: color_data = 12'h016;
			{9'd189, 8'd71}: color_data = 12'h027;
			{9'd189, 8'd72}: color_data = 12'h027;
			{9'd189, 8'd73}: color_data = 12'h027;
			{9'd189, 8'd74}: color_data = 12'h027;
			{9'd189, 8'd75}: color_data = 12'h028;
			{9'd189, 8'd76}: color_data = 12'h027;
			{9'd189, 8'd77}: color_data = 12'h001;
			{9'd189, 8'd119}: color_data = 12'h000;
			{9'd189, 8'd120}: color_data = 12'h016;
			{9'd189, 8'd121}: color_data = 12'h017;
			{9'd189, 8'd122}: color_data = 12'h017;
			{9'd189, 8'd123}: color_data = 12'h027;
			{9'd189, 8'd124}: color_data = 12'h027;
			{9'd189, 8'd125}: color_data = 12'h027;
			{9'd189, 8'd126}: color_data = 12'h027;
			{9'd189, 8'd127}: color_data = 12'h028;
			{9'd189, 8'd128}: color_data = 12'h014;
			{9'd189, 8'd129}: color_data = 12'h000;
			{9'd189, 8'd222}: color_data = 12'h300;
			{9'd189, 8'd223}: color_data = 12'hc30;
			{9'd189, 8'd224}: color_data = 12'hc30;
			{9'd189, 8'd225}: color_data = 12'h600;
			{9'd189, 8'd226}: color_data = 12'h100;
			{9'd189, 8'd227}: color_data = 12'h600;
			{9'd189, 8'd228}: color_data = 12'ha00;
			{9'd189, 8'd229}: color_data = 12'h900;
			{9'd189, 8'd230}: color_data = 12'h300;
			{9'd189, 8'd231}: color_data = 12'h620;
			{9'd189, 8'd232}: color_data = 12'hd40;
			{9'd189, 8'd233}: color_data = 12'ha20;
			{9'd189, 8'd234}: color_data = 12'h300;
			{9'd189, 8'd235}: color_data = 12'h200;
			{9'd189, 8'd236}: color_data = 12'h900;
			{9'd189, 8'd237}: color_data = 12'ha00;
			{9'd189, 8'd238}: color_data = 12'h700;
			{9'd189, 8'd239}: color_data = 12'h100;
			{9'd190, 8'd68}: color_data = 12'h035;
			{9'd190, 8'd69}: color_data = 12'h09e;
			{9'd190, 8'd70}: color_data = 12'h09e;
			{9'd190, 8'd71}: color_data = 12'h09e;
			{9'd190, 8'd72}: color_data = 12'h09e;
			{9'd190, 8'd73}: color_data = 12'h09e;
			{9'd190, 8'd74}: color_data = 12'h09e;
			{9'd190, 8'd75}: color_data = 12'h09e;
			{9'd190, 8'd76}: color_data = 12'h08c;
			{9'd190, 8'd77}: color_data = 12'h023;
			{9'd190, 8'd119}: color_data = 12'h000;
			{9'd190, 8'd120}: color_data = 12'h07b;
			{9'd190, 8'd121}: color_data = 12'h0ae;
			{9'd190, 8'd122}: color_data = 12'h09e;
			{9'd190, 8'd123}: color_data = 12'h09e;
			{9'd190, 8'd124}: color_data = 12'h09e;
			{9'd190, 8'd125}: color_data = 12'h09e;
			{9'd190, 8'd126}: color_data = 12'h09e;
			{9'd190, 8'd127}: color_data = 12'h09e;
			{9'd190, 8'd128}: color_data = 12'h057;
			{9'd190, 8'd129}: color_data = 12'h000;
			{9'd190, 8'd222}: color_data = 12'h000;
			{9'd190, 8'd223}: color_data = 12'h200;
			{9'd190, 8'd224}: color_data = 12'h300;
			{9'd190, 8'd225}: color_data = 12'h100;
			{9'd190, 8'd226}: color_data = 12'h000;
			{9'd190, 8'd227}: color_data = 12'h700;
			{9'd190, 8'd228}: color_data = 12'ha00;
			{9'd190, 8'd229}: color_data = 12'h900;
			{9'd190, 8'd230}: color_data = 12'h300;
			{9'd190, 8'd231}: color_data = 12'h100;
			{9'd190, 8'd232}: color_data = 12'h310;
			{9'd190, 8'd233}: color_data = 12'h200;
			{9'd190, 8'd234}: color_data = 12'h000;
			{9'd190, 8'd235}: color_data = 12'h300;
			{9'd190, 8'd236}: color_data = 12'h900;
			{9'd190, 8'd237}: color_data = 12'ha00;
			{9'd190, 8'd238}: color_data = 12'h700;
			{9'd190, 8'd239}: color_data = 12'h100;
			{9'd191, 8'd68}: color_data = 12'h057;
			{9'd191, 8'd69}: color_data = 12'h4ef;
			{9'd191, 8'd70}: color_data = 12'h7ef;
			{9'd191, 8'd71}: color_data = 12'h0cf;
			{9'd191, 8'd72}: color_data = 12'h0cf;
			{9'd191, 8'd73}: color_data = 12'h0df;
			{9'd191, 8'd74}: color_data = 12'h0bd;
			{9'd191, 8'd75}: color_data = 12'h068;
			{9'd191, 8'd76}: color_data = 12'h09c;
			{9'd191, 8'd77}: color_data = 12'h034;
			{9'd191, 8'd119}: color_data = 12'h000;
			{9'd191, 8'd120}: color_data = 12'h1ad;
			{9'd191, 8'd121}: color_data = 12'h8ff;
			{9'd191, 8'd122}: color_data = 12'h3df;
			{9'd191, 8'd123}: color_data = 12'h0cf;
			{9'd191, 8'd124}: color_data = 12'h0cf;
			{9'd191, 8'd125}: color_data = 12'h0cf;
			{9'd191, 8'd126}: color_data = 12'h07a;
			{9'd191, 8'd127}: color_data = 12'h08b;
			{9'd191, 8'd128}: color_data = 12'h079;
			{9'd191, 8'd129}: color_data = 12'h000;
			{9'd191, 8'd222}: color_data = 12'h100;
			{9'd191, 8'd223}: color_data = 12'h500;
			{9'd191, 8'd224}: color_data = 12'h500;
			{9'd191, 8'd225}: color_data = 12'h400;
			{9'd191, 8'd226}: color_data = 12'h100;
			{9'd191, 8'd227}: color_data = 12'ha20;
			{9'd191, 8'd228}: color_data = 12'hb10;
			{9'd191, 8'd229}: color_data = 12'h900;
			{9'd191, 8'd230}: color_data = 12'h300;
			{9'd191, 8'd231}: color_data = 12'h200;
			{9'd191, 8'd232}: color_data = 12'h500;
			{9'd191, 8'd233}: color_data = 12'h500;
			{9'd191, 8'd234}: color_data = 12'h200;
			{9'd191, 8'd235}: color_data = 12'h410;
			{9'd191, 8'd236}: color_data = 12'hc20;
			{9'd191, 8'd237}: color_data = 12'ha00;
			{9'd191, 8'd238}: color_data = 12'h700;
			{9'd191, 8'd239}: color_data = 12'h100;
			{9'd192, 8'd68}: color_data = 12'h047;
			{9'd192, 8'd69}: color_data = 12'h6df;
			{9'd192, 8'd70}: color_data = 12'heff;
			{9'd192, 8'd71}: color_data = 12'h6df;
			{9'd192, 8'd72}: color_data = 12'h0bf;
			{9'd192, 8'd73}: color_data = 12'h0bf;
			{9'd192, 8'd74}: color_data = 12'h056;
			{9'd192, 8'd75}: color_data = 12'h012;
			{9'd192, 8'd76}: color_data = 12'h08b;
			{9'd192, 8'd77}: color_data = 12'h034;
			{9'd192, 8'd119}: color_data = 12'h000;
			{9'd192, 8'd120}: color_data = 12'h2ac;
			{9'd192, 8'd121}: color_data = 12'hdff;
			{9'd192, 8'd122}: color_data = 12'haef;
			{9'd192, 8'd123}: color_data = 12'h1cf;
			{9'd192, 8'd124}: color_data = 12'h0cf;
			{9'd192, 8'd125}: color_data = 12'h08b;
			{9'd192, 8'd126}: color_data = 12'h012;
			{9'd192, 8'd127}: color_data = 12'h068;
			{9'd192, 8'd128}: color_data = 12'h079;
			{9'd192, 8'd129}: color_data = 12'h000;
			{9'd192, 8'd222}: color_data = 12'h200;
			{9'd192, 8'd223}: color_data = 12'h900;
			{9'd192, 8'd224}: color_data = 12'hb00;
			{9'd192, 8'd225}: color_data = 12'h800;
			{9'd192, 8'd226}: color_data = 12'h200;
			{9'd192, 8'd227}: color_data = 12'hb30;
			{9'd192, 8'd228}: color_data = 12'hc10;
			{9'd192, 8'd229}: color_data = 12'h800;
			{9'd192, 8'd230}: color_data = 12'h300;
			{9'd192, 8'd231}: color_data = 12'h400;
			{9'd192, 8'd232}: color_data = 12'ha00;
			{9'd192, 8'd233}: color_data = 12'ha00;
			{9'd192, 8'd234}: color_data = 12'h500;
			{9'd192, 8'd235}: color_data = 12'h510;
			{9'd192, 8'd236}: color_data = 12'hd30;
			{9'd192, 8'd237}: color_data = 12'ha00;
			{9'd192, 8'd238}: color_data = 12'h700;
			{9'd192, 8'd239}: color_data = 12'h100;
			{9'd193, 8'd68}: color_data = 12'h047;
			{9'd193, 8'd69}: color_data = 12'h6df;
			{9'd193, 8'd70}: color_data = 12'hfff;
			{9'd193, 8'd71}: color_data = 12'hdff;
			{9'd193, 8'd72}: color_data = 12'h5df;
			{9'd193, 8'd73}: color_data = 12'h068;
			{9'd193, 8'd74}: color_data = 12'h000;
			{9'd193, 8'd75}: color_data = 12'h012;
			{9'd193, 8'd76}: color_data = 12'h08c;
			{9'd193, 8'd77}: color_data = 12'h034;
			{9'd193, 8'd119}: color_data = 12'h000;
			{9'd193, 8'd120}: color_data = 12'h1ac;
			{9'd193, 8'd121}: color_data = 12'hdff;
			{9'd193, 8'd122}: color_data = 12'hfff;
			{9'd193, 8'd123}: color_data = 12'h9ef;
			{9'd193, 8'd124}: color_data = 12'h19c;
			{9'd193, 8'd125}: color_data = 12'h023;
			{9'd193, 8'd127}: color_data = 12'h068;
			{9'd193, 8'd128}: color_data = 12'h079;
			{9'd193, 8'd129}: color_data = 12'h000;
			{9'd193, 8'd222}: color_data = 12'h200;
			{9'd193, 8'd223}: color_data = 12'h900;
			{9'd193, 8'd224}: color_data = 12'ha00;
			{9'd193, 8'd225}: color_data = 12'h700;
			{9'd193, 8'd226}: color_data = 12'h200;
			{9'd193, 8'd227}: color_data = 12'hb30;
			{9'd193, 8'd228}: color_data = 12'he20;
			{9'd193, 8'd229}: color_data = 12'ha00;
			{9'd193, 8'd230}: color_data = 12'h300;
			{9'd193, 8'd231}: color_data = 12'h400;
			{9'd193, 8'd232}: color_data = 12'ha00;
			{9'd193, 8'd233}: color_data = 12'ha00;
			{9'd193, 8'd234}: color_data = 12'h400;
			{9'd193, 8'd235}: color_data = 12'h510;
			{9'd193, 8'd236}: color_data = 12'hf40;
			{9'd193, 8'd237}: color_data = 12'hd10;
			{9'd193, 8'd238}: color_data = 12'h800;
			{9'd193, 8'd239}: color_data = 12'h100;
			{9'd194, 8'd68}: color_data = 12'h047;
			{9'd194, 8'd69}: color_data = 12'h6df;
			{9'd194, 8'd70}: color_data = 12'hfff;
			{9'd194, 8'd71}: color_data = 12'hfff;
			{9'd194, 8'd72}: color_data = 12'h9aa;
			{9'd194, 8'd73}: color_data = 12'h011;
			{9'd194, 8'd75}: color_data = 12'h012;
			{9'd194, 8'd76}: color_data = 12'h08c;
			{9'd194, 8'd77}: color_data = 12'h034;
			{9'd194, 8'd119}: color_data = 12'h000;
			{9'd194, 8'd120}: color_data = 12'h1ac;
			{9'd194, 8'd121}: color_data = 12'hcff;
			{9'd194, 8'd122}: color_data = 12'hfff;
			{9'd194, 8'd123}: color_data = 12'hddd;
			{9'd194, 8'd124}: color_data = 12'h345;
			{9'd194, 8'd126}: color_data = 12'h000;
			{9'd194, 8'd127}: color_data = 12'h068;
			{9'd194, 8'd128}: color_data = 12'h079;
			{9'd194, 8'd129}: color_data = 12'h000;
			{9'd194, 8'd222}: color_data = 12'h200;
			{9'd194, 8'd223}: color_data = 12'h800;
			{9'd194, 8'd224}: color_data = 12'ha00;
			{9'd194, 8'd225}: color_data = 12'h800;
			{9'd194, 8'd226}: color_data = 12'h200;
			{9'd194, 8'd227}: color_data = 12'h930;
			{9'd194, 8'd228}: color_data = 12'hd30;
			{9'd194, 8'd229}: color_data = 12'h910;
			{9'd194, 8'd230}: color_data = 12'h200;
			{9'd194, 8'd231}: color_data = 12'h400;
			{9'd194, 8'd232}: color_data = 12'h900;
			{9'd194, 8'd233}: color_data = 12'ha00;
			{9'd194, 8'd234}: color_data = 12'h400;
			{9'd194, 8'd235}: color_data = 12'h310;
			{9'd194, 8'd236}: color_data = 12'hc30;
			{9'd194, 8'd237}: color_data = 12'hc20;
			{9'd194, 8'd238}: color_data = 12'h600;
			{9'd194, 8'd239}: color_data = 12'h000;
			{9'd195, 8'd68}: color_data = 12'h047;
			{9'd195, 8'd69}: color_data = 12'h6df;
			{9'd195, 8'd70}: color_data = 12'hfff;
			{9'd195, 8'd71}: color_data = 12'hcbb;
			{9'd195, 8'd72}: color_data = 12'h323;
			{9'd195, 8'd73}: color_data = 12'h002;
			{9'd195, 8'd74}: color_data = 12'h000;
			{9'd195, 8'd75}: color_data = 12'h012;
			{9'd195, 8'd76}: color_data = 12'h08c;
			{9'd195, 8'd77}: color_data = 12'h034;
			{9'd195, 8'd119}: color_data = 12'h000;
			{9'd195, 8'd120}: color_data = 12'h1ac;
			{9'd195, 8'd121}: color_data = 12'hdff;
			{9'd195, 8'd122}: color_data = 12'hfee;
			{9'd195, 8'd123}: color_data = 12'h666;
			{9'd195, 8'd124}: color_data = 12'h002;
			{9'd195, 8'd125}: color_data = 12'h001;
			{9'd195, 8'd126}: color_data = 12'h000;
			{9'd195, 8'd127}: color_data = 12'h068;
			{9'd195, 8'd128}: color_data = 12'h079;
			{9'd195, 8'd129}: color_data = 12'h000;
			{9'd195, 8'd222}: color_data = 12'h200;
			{9'd195, 8'd223}: color_data = 12'h900;
			{9'd195, 8'd224}: color_data = 12'ha00;
			{9'd195, 8'd225}: color_data = 12'h800;
			{9'd195, 8'd226}: color_data = 12'h100;
			{9'd195, 8'd227}: color_data = 12'h100;
			{9'd195, 8'd228}: color_data = 12'h310;
			{9'd195, 8'd229}: color_data = 12'h200;
			{9'd195, 8'd230}: color_data = 12'h000;
			{9'd195, 8'd231}: color_data = 12'h500;
			{9'd195, 8'd232}: color_data = 12'ha00;
			{9'd195, 8'd233}: color_data = 12'ha00;
			{9'd195, 8'd234}: color_data = 12'h500;
			{9'd195, 8'd235}: color_data = 12'h000;
			{9'd195, 8'd236}: color_data = 12'h200;
			{9'd195, 8'd237}: color_data = 12'h300;
			{9'd195, 8'd238}: color_data = 12'h100;
			{9'd195, 8'd239}: color_data = 12'h000;
			{9'd196, 8'd68}: color_data = 12'h047;
			{9'd196, 8'd69}: color_data = 12'h6ef;
			{9'd196, 8'd70}: color_data = 12'hdcc;
			{9'd196, 8'd71}: color_data = 12'h434;
			{9'd196, 8'd72}: color_data = 12'h003;
			{9'd196, 8'd73}: color_data = 12'h005;
			{9'd196, 8'd74}: color_data = 12'h002;
			{9'd196, 8'd75}: color_data = 12'h012;
			{9'd196, 8'd76}: color_data = 12'h08c;
			{9'd196, 8'd77}: color_data = 12'h034;
			{9'd196, 8'd119}: color_data = 12'h000;
			{9'd196, 8'd120}: color_data = 12'h2ad;
			{9'd196, 8'd121}: color_data = 12'hcff;
			{9'd196, 8'd122}: color_data = 12'h877;
			{9'd196, 8'd123}: color_data = 12'h002;
			{9'd196, 8'd124}: color_data = 12'h004;
			{9'd196, 8'd125}: color_data = 12'h004;
			{9'd196, 8'd126}: color_data = 12'h000;
			{9'd196, 8'd127}: color_data = 12'h068;
			{9'd196, 8'd128}: color_data = 12'h079;
			{9'd196, 8'd129}: color_data = 12'h000;
			{9'd196, 8'd222}: color_data = 12'h300;
			{9'd196, 8'd223}: color_data = 12'hc20;
			{9'd196, 8'd224}: color_data = 12'ha00;
			{9'd196, 8'd225}: color_data = 12'h800;
			{9'd196, 8'd226}: color_data = 12'h100;
			{9'd196, 8'd227}: color_data = 12'h300;
			{9'd196, 8'd228}: color_data = 12'h500;
			{9'd196, 8'd229}: color_data = 12'h500;
			{9'd196, 8'd230}: color_data = 12'h100;
			{9'd196, 8'd231}: color_data = 12'h710;
			{9'd196, 8'd232}: color_data = 12'hc10;
			{9'd196, 8'd233}: color_data = 12'h900;
			{9'd196, 8'd234}: color_data = 12'h500;
			{9'd196, 8'd235}: color_data = 12'h100;
			{9'd196, 8'd236}: color_data = 12'h500;
			{9'd196, 8'd237}: color_data = 12'h600;
			{9'd196, 8'd238}: color_data = 12'h400;
			{9'd196, 8'd239}: color_data = 12'h000;
			{9'd197, 8'd68}: color_data = 12'h057;
			{9'd197, 8'd69}: color_data = 12'h3bd;
			{9'd197, 8'd70}: color_data = 12'h555;
			{9'd197, 8'd71}: color_data = 12'h002;
			{9'd197, 8'd72}: color_data = 12'h005;
			{9'd197, 8'd73}: color_data = 12'h005;
			{9'd197, 8'd74}: color_data = 12'h004;
			{9'd197, 8'd75}: color_data = 12'h025;
			{9'd197, 8'd76}: color_data = 12'h09c;
			{9'd197, 8'd77}: color_data = 12'h034;
			{9'd197, 8'd119}: color_data = 12'h000;
			{9'd197, 8'd120}: color_data = 12'h1ac;
			{9'd197, 8'd121}: color_data = 12'h689;
			{9'd197, 8'd122}: color_data = 12'h212;
			{9'd197, 8'd123}: color_data = 12'h004;
			{9'd197, 8'd124}: color_data = 12'h005;
			{9'd197, 8'd125}: color_data = 12'h005;
			{9'd197, 8'd126}: color_data = 12'h003;
			{9'd197, 8'd127}: color_data = 12'h06a;
			{9'd197, 8'd128}: color_data = 12'h079;
			{9'd197, 8'd129}: color_data = 12'h000;
			{9'd197, 8'd222}: color_data = 12'h410;
			{9'd197, 8'd223}: color_data = 12'hd30;
			{9'd197, 8'd224}: color_data = 12'hb00;
			{9'd197, 8'd225}: color_data = 12'h700;
			{9'd197, 8'd226}: color_data = 12'h200;
			{9'd197, 8'd227}: color_data = 12'h700;
			{9'd197, 8'd228}: color_data = 12'hb00;
			{9'd197, 8'd229}: color_data = 12'h900;
			{9'd197, 8'd230}: color_data = 12'h300;
			{9'd197, 8'd231}: color_data = 12'h820;
			{9'd197, 8'd232}: color_data = 12'hd20;
			{9'd197, 8'd233}: color_data = 12'h900;
			{9'd197, 8'd234}: color_data = 12'h500;
			{9'd197, 8'd235}: color_data = 12'h300;
			{9'd197, 8'd236}: color_data = 12'h900;
			{9'd197, 8'd237}: color_data = 12'hb00;
			{9'd197, 8'd238}: color_data = 12'h800;
			{9'd197, 8'd239}: color_data = 12'h100;
			{9'd198, 8'd68}: color_data = 12'h035;
			{9'd198, 8'd69}: color_data = 12'h047;
			{9'd198, 8'd70}: color_data = 12'h001;
			{9'd198, 8'd71}: color_data = 12'h004;
			{9'd198, 8'd72}: color_data = 12'h004;
			{9'd198, 8'd73}: color_data = 12'h004;
			{9'd198, 8'd74}: color_data = 12'h004;
			{9'd198, 8'd75}: color_data = 12'h015;
			{9'd198, 8'd76}: color_data = 12'h059;
			{9'd198, 8'd77}: color_data = 12'h023;
			{9'd198, 8'd119}: color_data = 12'h000;
			{9'd198, 8'd120}: color_data = 12'h048;
			{9'd198, 8'd121}: color_data = 12'h013;
			{9'd198, 8'd122}: color_data = 12'h002;
			{9'd198, 8'd123}: color_data = 12'h004;
			{9'd198, 8'd124}: color_data = 12'h004;
			{9'd198, 8'd125}: color_data = 12'h004;
			{9'd198, 8'd126}: color_data = 12'h004;
			{9'd198, 8'd127}: color_data = 12'h038;
			{9'd198, 8'd128}: color_data = 12'h046;
			{9'd198, 8'd129}: color_data = 12'h000;
			{9'd198, 8'd222}: color_data = 12'h410;
			{9'd198, 8'd223}: color_data = 12'he40;
			{9'd198, 8'd224}: color_data = 12'hd20;
			{9'd198, 8'd225}: color_data = 12'h800;
			{9'd198, 8'd226}: color_data = 12'h200;
			{9'd198, 8'd227}: color_data = 12'h600;
			{9'd198, 8'd228}: color_data = 12'ha00;
			{9'd198, 8'd229}: color_data = 12'h900;
			{9'd198, 8'd230}: color_data = 12'h300;
			{9'd198, 8'd231}: color_data = 12'h820;
			{9'd198, 8'd232}: color_data = 12'hf30;
			{9'd198, 8'd233}: color_data = 12'hc00;
			{9'd198, 8'd234}: color_data = 12'h500;
			{9'd198, 8'd235}: color_data = 12'h200;
			{9'd198, 8'd236}: color_data = 12'h900;
			{9'd198, 8'd237}: color_data = 12'ha00;
			{9'd198, 8'd238}: color_data = 12'h700;
			{9'd198, 8'd239}: color_data = 12'h100;
			{9'd199, 8'd68}: color_data = 12'h013;
			{9'd199, 8'd69}: color_data = 12'h027;
			{9'd199, 8'd70}: color_data = 12'h016;
			{9'd199, 8'd71}: color_data = 12'h027;
			{9'd199, 8'd72}: color_data = 12'h027;
			{9'd199, 8'd73}: color_data = 12'h027;
			{9'd199, 8'd74}: color_data = 12'h027;
			{9'd199, 8'd75}: color_data = 12'h028;
			{9'd199, 8'd76}: color_data = 12'h027;
			{9'd199, 8'd77}: color_data = 12'h001;
			{9'd199, 8'd119}: color_data = 12'h000;
			{9'd199, 8'd120}: color_data = 12'h015;
			{9'd199, 8'd121}: color_data = 12'h027;
			{9'd199, 8'd122}: color_data = 12'h026;
			{9'd199, 8'd123}: color_data = 12'h027;
			{9'd199, 8'd124}: color_data = 12'h027;
			{9'd199, 8'd125}: color_data = 12'h027;
			{9'd199, 8'd126}: color_data = 12'h027;
			{9'd199, 8'd127}: color_data = 12'h028;
			{9'd199, 8'd128}: color_data = 12'h014;
			{9'd199, 8'd129}: color_data = 12'h000;
			{9'd199, 8'd222}: color_data = 12'h300;
			{9'd199, 8'd223}: color_data = 12'hc30;
			{9'd199, 8'd224}: color_data = 12'hc30;
			{9'd199, 8'd225}: color_data = 12'h600;
			{9'd199, 8'd226}: color_data = 12'h100;
			{9'd199, 8'd227}: color_data = 12'h600;
			{9'd199, 8'd228}: color_data = 12'ha00;
			{9'd199, 8'd229}: color_data = 12'h900;
			{9'd199, 8'd230}: color_data = 12'h300;
			{9'd199, 8'd231}: color_data = 12'h620;
			{9'd199, 8'd232}: color_data = 12'hd40;
			{9'd199, 8'd233}: color_data = 12'ha20;
			{9'd199, 8'd234}: color_data = 12'h300;
			{9'd199, 8'd235}: color_data = 12'h200;
			{9'd199, 8'd236}: color_data = 12'h900;
			{9'd199, 8'd237}: color_data = 12'ha00;
			{9'd199, 8'd238}: color_data = 12'h700;
			{9'd199, 8'd239}: color_data = 12'h100;
			{9'd200, 8'd68}: color_data = 12'h036;
			{9'd200, 8'd69}: color_data = 12'h09e;
			{9'd200, 8'd70}: color_data = 12'h09e;
			{9'd200, 8'd71}: color_data = 12'h09e;
			{9'd200, 8'd72}: color_data = 12'h09e;
			{9'd200, 8'd73}: color_data = 12'h09e;
			{9'd200, 8'd74}: color_data = 12'h09e;
			{9'd200, 8'd75}: color_data = 12'h09e;
			{9'd200, 8'd76}: color_data = 12'h08c;
			{9'd200, 8'd77}: color_data = 12'h023;
			{9'd200, 8'd119}: color_data = 12'h000;
			{9'd200, 8'd120}: color_data = 12'h07b;
			{9'd200, 8'd121}: color_data = 12'h0ae;
			{9'd200, 8'd122}: color_data = 12'h09e;
			{9'd200, 8'd123}: color_data = 12'h09e;
			{9'd200, 8'd124}: color_data = 12'h09e;
			{9'd200, 8'd125}: color_data = 12'h09e;
			{9'd200, 8'd126}: color_data = 12'h09e;
			{9'd200, 8'd127}: color_data = 12'h09e;
			{9'd200, 8'd128}: color_data = 12'h057;
			{9'd200, 8'd129}: color_data = 12'h000;
			{9'd200, 8'd222}: color_data = 12'h000;
			{9'd200, 8'd223}: color_data = 12'h200;
			{9'd200, 8'd224}: color_data = 12'h300;
			{9'd200, 8'd225}: color_data = 12'h100;
			{9'd200, 8'd226}: color_data = 12'h000;
			{9'd200, 8'd227}: color_data = 12'h700;
			{9'd200, 8'd228}: color_data = 12'ha00;
			{9'd200, 8'd229}: color_data = 12'h900;
			{9'd200, 8'd230}: color_data = 12'h300;
			{9'd200, 8'd231}: color_data = 12'h000;
			{9'd200, 8'd232}: color_data = 12'h300;
			{9'd200, 8'd233}: color_data = 12'h200;
			{9'd200, 8'd234}: color_data = 12'h000;
			{9'd200, 8'd235}: color_data = 12'h300;
			{9'd200, 8'd236}: color_data = 12'h900;
			{9'd200, 8'd237}: color_data = 12'ha00;
			{9'd200, 8'd238}: color_data = 12'h700;
			{9'd200, 8'd239}: color_data = 12'h100;
			{9'd201, 8'd68}: color_data = 12'h057;
			{9'd201, 8'd69}: color_data = 12'h4ef;
			{9'd201, 8'd70}: color_data = 12'h7ef;
			{9'd201, 8'd71}: color_data = 12'h0cf;
			{9'd201, 8'd72}: color_data = 12'h0cf;
			{9'd201, 8'd73}: color_data = 12'h0df;
			{9'd201, 8'd74}: color_data = 12'h0bd;
			{9'd201, 8'd75}: color_data = 12'h068;
			{9'd201, 8'd76}: color_data = 12'h09c;
			{9'd201, 8'd77}: color_data = 12'h034;
			{9'd201, 8'd119}: color_data = 12'h000;
			{9'd201, 8'd120}: color_data = 12'h1ad;
			{9'd201, 8'd121}: color_data = 12'h8ff;
			{9'd201, 8'd122}: color_data = 12'h3df;
			{9'd201, 8'd123}: color_data = 12'h0cf;
			{9'd201, 8'd124}: color_data = 12'h0cf;
			{9'd201, 8'd125}: color_data = 12'h0cf;
			{9'd201, 8'd126}: color_data = 12'h079;
			{9'd201, 8'd127}: color_data = 12'h08b;
			{9'd201, 8'd128}: color_data = 12'h079;
			{9'd201, 8'd129}: color_data = 12'h000;
			{9'd201, 8'd222}: color_data = 12'h100;
			{9'd201, 8'd223}: color_data = 12'h500;
			{9'd201, 8'd224}: color_data = 12'h600;
			{9'd201, 8'd225}: color_data = 12'h400;
			{9'd201, 8'd226}: color_data = 12'h200;
			{9'd201, 8'd227}: color_data = 12'ha20;
			{9'd201, 8'd228}: color_data = 12'hb10;
			{9'd201, 8'd229}: color_data = 12'h900;
			{9'd201, 8'd230}: color_data = 12'h300;
			{9'd201, 8'd231}: color_data = 12'h200;
			{9'd201, 8'd232}: color_data = 12'h500;
			{9'd201, 8'd233}: color_data = 12'h500;
			{9'd201, 8'd234}: color_data = 12'h200;
			{9'd201, 8'd235}: color_data = 12'h410;
			{9'd201, 8'd236}: color_data = 12'hc20;
			{9'd201, 8'd237}: color_data = 12'ha00;
			{9'd201, 8'd238}: color_data = 12'h700;
			{9'd201, 8'd239}: color_data = 12'h100;
			{9'd202, 8'd68}: color_data = 12'h047;
			{9'd202, 8'd69}: color_data = 12'h6df;
			{9'd202, 8'd70}: color_data = 12'heff;
			{9'd202, 8'd71}: color_data = 12'h6df;
			{9'd202, 8'd72}: color_data = 12'h0bf;
			{9'd202, 8'd73}: color_data = 12'h0bf;
			{9'd202, 8'd74}: color_data = 12'h056;
			{9'd202, 8'd75}: color_data = 12'h012;
			{9'd202, 8'd76}: color_data = 12'h08b;
			{9'd202, 8'd77}: color_data = 12'h034;
			{9'd202, 8'd119}: color_data = 12'h000;
			{9'd202, 8'd120}: color_data = 12'h2ac;
			{9'd202, 8'd121}: color_data = 12'hdff;
			{9'd202, 8'd122}: color_data = 12'haef;
			{9'd202, 8'd123}: color_data = 12'h1cf;
			{9'd202, 8'd124}: color_data = 12'h0cf;
			{9'd202, 8'd125}: color_data = 12'h08b;
			{9'd202, 8'd126}: color_data = 12'h012;
			{9'd202, 8'd127}: color_data = 12'h068;
			{9'd202, 8'd128}: color_data = 12'h079;
			{9'd202, 8'd129}: color_data = 12'h000;
			{9'd202, 8'd222}: color_data = 12'h200;
			{9'd202, 8'd223}: color_data = 12'h900;
			{9'd202, 8'd224}: color_data = 12'hb00;
			{9'd202, 8'd225}: color_data = 12'h800;
			{9'd202, 8'd226}: color_data = 12'h200;
			{9'd202, 8'd227}: color_data = 12'hb30;
			{9'd202, 8'd228}: color_data = 12'hc10;
			{9'd202, 8'd229}: color_data = 12'h800;
			{9'd202, 8'd230}: color_data = 12'h300;
			{9'd202, 8'd231}: color_data = 12'h400;
			{9'd202, 8'd232}: color_data = 12'ha00;
			{9'd202, 8'd233}: color_data = 12'ha00;
			{9'd202, 8'd234}: color_data = 12'h500;
			{9'd202, 8'd235}: color_data = 12'h510;
			{9'd202, 8'd236}: color_data = 12'hd30;
			{9'd202, 8'd237}: color_data = 12'ha00;
			{9'd202, 8'd238}: color_data = 12'h700;
			{9'd202, 8'd239}: color_data = 12'h100;
			{9'd203, 8'd68}: color_data = 12'h047;
			{9'd203, 8'd69}: color_data = 12'h6df;
			{9'd203, 8'd70}: color_data = 12'hfff;
			{9'd203, 8'd71}: color_data = 12'hdff;
			{9'd203, 8'd72}: color_data = 12'h5df;
			{9'd203, 8'd73}: color_data = 12'h068;
			{9'd203, 8'd74}: color_data = 12'h000;
			{9'd203, 8'd75}: color_data = 12'h012;
			{9'd203, 8'd76}: color_data = 12'h08c;
			{9'd203, 8'd77}: color_data = 12'h034;
			{9'd203, 8'd119}: color_data = 12'h000;
			{9'd203, 8'd120}: color_data = 12'h1ac;
			{9'd203, 8'd121}: color_data = 12'hdff;
			{9'd203, 8'd122}: color_data = 12'hfff;
			{9'd203, 8'd123}: color_data = 12'h8ef;
			{9'd203, 8'd124}: color_data = 12'h19c;
			{9'd203, 8'd125}: color_data = 12'h023;
			{9'd203, 8'd127}: color_data = 12'h068;
			{9'd203, 8'd128}: color_data = 12'h079;
			{9'd203, 8'd129}: color_data = 12'h000;
			{9'd203, 8'd222}: color_data = 12'h200;
			{9'd203, 8'd223}: color_data = 12'h900;
			{9'd203, 8'd224}: color_data = 12'ha00;
			{9'd203, 8'd225}: color_data = 12'h700;
			{9'd203, 8'd226}: color_data = 12'h200;
			{9'd203, 8'd227}: color_data = 12'hb30;
			{9'd203, 8'd228}: color_data = 12'he20;
			{9'd203, 8'd229}: color_data = 12'ha00;
			{9'd203, 8'd230}: color_data = 12'h300;
			{9'd203, 8'd231}: color_data = 12'h400;
			{9'd203, 8'd232}: color_data = 12'ha00;
			{9'd203, 8'd233}: color_data = 12'ha00;
			{9'd203, 8'd234}: color_data = 12'h400;
			{9'd203, 8'd235}: color_data = 12'h510;
			{9'd203, 8'd236}: color_data = 12'hf40;
			{9'd203, 8'd237}: color_data = 12'hd10;
			{9'd203, 8'd238}: color_data = 12'h800;
			{9'd203, 8'd239}: color_data = 12'h100;
			{9'd204, 8'd68}: color_data = 12'h047;
			{9'd204, 8'd69}: color_data = 12'h6df;
			{9'd204, 8'd70}: color_data = 12'hfff;
			{9'd204, 8'd71}: color_data = 12'hfff;
			{9'd204, 8'd72}: color_data = 12'h9aa;
			{9'd204, 8'd73}: color_data = 12'h011;
			{9'd204, 8'd75}: color_data = 12'h012;
			{9'd204, 8'd76}: color_data = 12'h08c;
			{9'd204, 8'd77}: color_data = 12'h034;
			{9'd204, 8'd119}: color_data = 12'h000;
			{9'd204, 8'd120}: color_data = 12'h1ac;
			{9'd204, 8'd121}: color_data = 12'hcff;
			{9'd204, 8'd122}: color_data = 12'hfff;
			{9'd204, 8'd123}: color_data = 12'hddd;
			{9'd204, 8'd124}: color_data = 12'h345;
			{9'd204, 8'd126}: color_data = 12'h000;
			{9'd204, 8'd127}: color_data = 12'h068;
			{9'd204, 8'd128}: color_data = 12'h079;
			{9'd204, 8'd129}: color_data = 12'h000;
			{9'd204, 8'd222}: color_data = 12'h200;
			{9'd204, 8'd223}: color_data = 12'h800;
			{9'd204, 8'd224}: color_data = 12'ha00;
			{9'd204, 8'd225}: color_data = 12'h800;
			{9'd204, 8'd226}: color_data = 12'h200;
			{9'd204, 8'd227}: color_data = 12'h920;
			{9'd204, 8'd228}: color_data = 12'hd30;
			{9'd204, 8'd229}: color_data = 12'h910;
			{9'd204, 8'd230}: color_data = 12'h200;
			{9'd204, 8'd231}: color_data = 12'h400;
			{9'd204, 8'd232}: color_data = 12'h900;
			{9'd204, 8'd233}: color_data = 12'ha00;
			{9'd204, 8'd234}: color_data = 12'h400;
			{9'd204, 8'd235}: color_data = 12'h310;
			{9'd204, 8'd236}: color_data = 12'hc30;
			{9'd204, 8'd237}: color_data = 12'hc20;
			{9'd204, 8'd238}: color_data = 12'h600;
			{9'd204, 8'd239}: color_data = 12'h000;
			{9'd205, 8'd68}: color_data = 12'h047;
			{9'd205, 8'd69}: color_data = 12'h6df;
			{9'd205, 8'd70}: color_data = 12'hfff;
			{9'd205, 8'd71}: color_data = 12'hcbb;
			{9'd205, 8'd72}: color_data = 12'h323;
			{9'd205, 8'd73}: color_data = 12'h002;
			{9'd205, 8'd74}: color_data = 12'h000;
			{9'd205, 8'd75}: color_data = 12'h012;
			{9'd205, 8'd76}: color_data = 12'h08c;
			{9'd205, 8'd77}: color_data = 12'h034;
			{9'd205, 8'd119}: color_data = 12'h000;
			{9'd205, 8'd120}: color_data = 12'h1ac;
			{9'd205, 8'd121}: color_data = 12'hdff;
			{9'd205, 8'd122}: color_data = 12'hfee;
			{9'd205, 8'd123}: color_data = 12'h666;
			{9'd205, 8'd124}: color_data = 12'h002;
			{9'd205, 8'd125}: color_data = 12'h001;
			{9'd205, 8'd126}: color_data = 12'h000;
			{9'd205, 8'd127}: color_data = 12'h068;
			{9'd205, 8'd128}: color_data = 12'h079;
			{9'd205, 8'd129}: color_data = 12'h000;
			{9'd205, 8'd222}: color_data = 12'h200;
			{9'd205, 8'd223}: color_data = 12'h900;
			{9'd205, 8'd224}: color_data = 12'ha00;
			{9'd205, 8'd225}: color_data = 12'h800;
			{9'd205, 8'd226}: color_data = 12'h100;
			{9'd205, 8'd227}: color_data = 12'h100;
			{9'd205, 8'd228}: color_data = 12'h310;
			{9'd205, 8'd229}: color_data = 12'h200;
			{9'd205, 8'd230}: color_data = 12'h000;
			{9'd205, 8'd231}: color_data = 12'h500;
			{9'd205, 8'd232}: color_data = 12'ha00;
			{9'd205, 8'd233}: color_data = 12'ha00;
			{9'd205, 8'd234}: color_data = 12'h500;
			{9'd205, 8'd235}: color_data = 12'h000;
			{9'd205, 8'd236}: color_data = 12'h200;
			{9'd205, 8'd237}: color_data = 12'h300;
			{9'd205, 8'd238}: color_data = 12'h100;
			{9'd205, 8'd239}: color_data = 12'h000;
			{9'd206, 8'd68}: color_data = 12'h047;
			{9'd206, 8'd69}: color_data = 12'h6ef;
			{9'd206, 8'd70}: color_data = 12'hddc;
			{9'd206, 8'd71}: color_data = 12'h434;
			{9'd206, 8'd72}: color_data = 12'h003;
			{9'd206, 8'd73}: color_data = 12'h005;
			{9'd206, 8'd74}: color_data = 12'h002;
			{9'd206, 8'd75}: color_data = 12'h012;
			{9'd206, 8'd76}: color_data = 12'h08c;
			{9'd206, 8'd77}: color_data = 12'h034;
			{9'd206, 8'd119}: color_data = 12'h000;
			{9'd206, 8'd120}: color_data = 12'h2ad;
			{9'd206, 8'd121}: color_data = 12'hcff;
			{9'd206, 8'd122}: color_data = 12'h877;
			{9'd206, 8'd123}: color_data = 12'h002;
			{9'd206, 8'd124}: color_data = 12'h004;
			{9'd206, 8'd125}: color_data = 12'h004;
			{9'd206, 8'd126}: color_data = 12'h000;
			{9'd206, 8'd127}: color_data = 12'h068;
			{9'd206, 8'd128}: color_data = 12'h079;
			{9'd206, 8'd129}: color_data = 12'h000;
			{9'd206, 8'd222}: color_data = 12'h300;
			{9'd206, 8'd223}: color_data = 12'hc20;
			{9'd206, 8'd224}: color_data = 12'ha00;
			{9'd206, 8'd225}: color_data = 12'h800;
			{9'd206, 8'd226}: color_data = 12'h100;
			{9'd206, 8'd227}: color_data = 12'h300;
			{9'd206, 8'd228}: color_data = 12'h500;
			{9'd206, 8'd229}: color_data = 12'h500;
			{9'd206, 8'd230}: color_data = 12'h100;
			{9'd206, 8'd231}: color_data = 12'h710;
			{9'd206, 8'd232}: color_data = 12'hc10;
			{9'd206, 8'd233}: color_data = 12'h900;
			{9'd206, 8'd234}: color_data = 12'h500;
			{9'd206, 8'd235}: color_data = 12'h100;
			{9'd206, 8'd236}: color_data = 12'h500;
			{9'd206, 8'd237}: color_data = 12'h600;
			{9'd206, 8'd238}: color_data = 12'h400;
			{9'd206, 8'd239}: color_data = 12'h000;
			{9'd207, 8'd68}: color_data = 12'h057;
			{9'd207, 8'd69}: color_data = 12'h3bd;
			{9'd207, 8'd70}: color_data = 12'h555;
			{9'd207, 8'd71}: color_data = 12'h002;
			{9'd207, 8'd72}: color_data = 12'h005;
			{9'd207, 8'd73}: color_data = 12'h005;
			{9'd207, 8'd74}: color_data = 12'h004;
			{9'd207, 8'd75}: color_data = 12'h025;
			{9'd207, 8'd76}: color_data = 12'h09c;
			{9'd207, 8'd77}: color_data = 12'h034;
			{9'd207, 8'd119}: color_data = 12'h000;
			{9'd207, 8'd120}: color_data = 12'h1ac;
			{9'd207, 8'd121}: color_data = 12'h689;
			{9'd207, 8'd122}: color_data = 12'h212;
			{9'd207, 8'd123}: color_data = 12'h004;
			{9'd207, 8'd124}: color_data = 12'h005;
			{9'd207, 8'd125}: color_data = 12'h005;
			{9'd207, 8'd126}: color_data = 12'h003;
			{9'd207, 8'd127}: color_data = 12'h06a;
			{9'd207, 8'd128}: color_data = 12'h079;
			{9'd207, 8'd129}: color_data = 12'h000;
			{9'd207, 8'd222}: color_data = 12'h410;
			{9'd207, 8'd223}: color_data = 12'hd30;
			{9'd207, 8'd224}: color_data = 12'hb00;
			{9'd207, 8'd225}: color_data = 12'h700;
			{9'd207, 8'd226}: color_data = 12'h200;
			{9'd207, 8'd227}: color_data = 12'h700;
			{9'd207, 8'd228}: color_data = 12'hb00;
			{9'd207, 8'd229}: color_data = 12'ha00;
			{9'd207, 8'd230}: color_data = 12'h300;
			{9'd207, 8'd231}: color_data = 12'h820;
			{9'd207, 8'd232}: color_data = 12'hd20;
			{9'd207, 8'd233}: color_data = 12'h900;
			{9'd207, 8'd234}: color_data = 12'h500;
			{9'd207, 8'd235}: color_data = 12'h300;
			{9'd207, 8'd236}: color_data = 12'h900;
			{9'd207, 8'd237}: color_data = 12'hb00;
			{9'd207, 8'd238}: color_data = 12'h800;
			{9'd207, 8'd239}: color_data = 12'h100;
			{9'd208, 8'd68}: color_data = 12'h035;
			{9'd208, 8'd69}: color_data = 12'h047;
			{9'd208, 8'd70}: color_data = 12'h001;
			{9'd208, 8'd71}: color_data = 12'h004;
			{9'd208, 8'd72}: color_data = 12'h004;
			{9'd208, 8'd73}: color_data = 12'h004;
			{9'd208, 8'd74}: color_data = 12'h004;
			{9'd208, 8'd75}: color_data = 12'h015;
			{9'd208, 8'd76}: color_data = 12'h059;
			{9'd208, 8'd77}: color_data = 12'h023;
			{9'd208, 8'd119}: color_data = 12'h000;
			{9'd208, 8'd120}: color_data = 12'h058;
			{9'd208, 8'd121}: color_data = 12'h013;
			{9'd208, 8'd122}: color_data = 12'h002;
			{9'd208, 8'd123}: color_data = 12'h004;
			{9'd208, 8'd124}: color_data = 12'h004;
			{9'd208, 8'd125}: color_data = 12'h004;
			{9'd208, 8'd126}: color_data = 12'h004;
			{9'd208, 8'd127}: color_data = 12'h039;
			{9'd208, 8'd128}: color_data = 12'h046;
			{9'd208, 8'd129}: color_data = 12'h000;
			{9'd208, 8'd222}: color_data = 12'h410;
			{9'd208, 8'd223}: color_data = 12'he40;
			{9'd208, 8'd224}: color_data = 12'hd20;
			{9'd208, 8'd225}: color_data = 12'h800;
			{9'd208, 8'd226}: color_data = 12'h200;
			{9'd208, 8'd227}: color_data = 12'h600;
			{9'd208, 8'd228}: color_data = 12'ha00;
			{9'd208, 8'd229}: color_data = 12'h900;
			{9'd208, 8'd230}: color_data = 12'h300;
			{9'd208, 8'd231}: color_data = 12'h820;
			{9'd208, 8'd232}: color_data = 12'hf30;
			{9'd208, 8'd233}: color_data = 12'hc00;
			{9'd208, 8'd234}: color_data = 12'h500;
			{9'd208, 8'd235}: color_data = 12'h200;
			{9'd208, 8'd236}: color_data = 12'h900;
			{9'd208, 8'd237}: color_data = 12'ha00;
			{9'd208, 8'd238}: color_data = 12'h700;
			{9'd208, 8'd239}: color_data = 12'h100;
			{9'd209, 8'd68}: color_data = 12'h013;
			{9'd209, 8'd69}: color_data = 12'h027;
			{9'd209, 8'd70}: color_data = 12'h016;
			{9'd209, 8'd71}: color_data = 12'h027;
			{9'd209, 8'd72}: color_data = 12'h027;
			{9'd209, 8'd73}: color_data = 12'h017;
			{9'd209, 8'd74}: color_data = 12'h027;
			{9'd209, 8'd75}: color_data = 12'h028;
			{9'd209, 8'd76}: color_data = 12'h027;
			{9'd209, 8'd77}: color_data = 12'h001;
			{9'd209, 8'd119}: color_data = 12'h000;
			{9'd209, 8'd120}: color_data = 12'h016;
			{9'd209, 8'd121}: color_data = 12'h017;
			{9'd209, 8'd122}: color_data = 12'h016;
			{9'd209, 8'd123}: color_data = 12'h027;
			{9'd209, 8'd124}: color_data = 12'h027;
			{9'd209, 8'd125}: color_data = 12'h017;
			{9'd209, 8'd126}: color_data = 12'h027;
			{9'd209, 8'd127}: color_data = 12'h028;
			{9'd209, 8'd128}: color_data = 12'h014;
			{9'd209, 8'd129}: color_data = 12'h000;
			{9'd209, 8'd171}: color_data = 12'h011;
			{9'd209, 8'd172}: color_data = 12'h023;
			{9'd209, 8'd173}: color_data = 12'h012;
			{9'd209, 8'd174}: color_data = 12'h022;
			{9'd209, 8'd175}: color_data = 12'h022;
			{9'd209, 8'd176}: color_data = 12'h012;
			{9'd209, 8'd177}: color_data = 12'h023;
			{9'd209, 8'd178}: color_data = 12'h023;
			{9'd209, 8'd179}: color_data = 12'h012;
			{9'd209, 8'd180}: color_data = 12'h000;
			{9'd209, 8'd222}: color_data = 12'h300;
			{9'd209, 8'd223}: color_data = 12'hc30;
			{9'd209, 8'd224}: color_data = 12'hc30;
			{9'd209, 8'd225}: color_data = 12'h600;
			{9'd209, 8'd226}: color_data = 12'h100;
			{9'd209, 8'd227}: color_data = 12'h600;
			{9'd209, 8'd228}: color_data = 12'ha00;
			{9'd209, 8'd229}: color_data = 12'h900;
			{9'd209, 8'd230}: color_data = 12'h300;
			{9'd209, 8'd231}: color_data = 12'h620;
			{9'd209, 8'd232}: color_data = 12'hd40;
			{9'd209, 8'd233}: color_data = 12'ha20;
			{9'd209, 8'd234}: color_data = 12'h300;
			{9'd209, 8'd235}: color_data = 12'h200;
			{9'd209, 8'd236}: color_data = 12'h900;
			{9'd209, 8'd237}: color_data = 12'ha00;
			{9'd209, 8'd238}: color_data = 12'h700;
			{9'd209, 8'd239}: color_data = 12'h100;
			{9'd210, 8'd68}: color_data = 12'h045;
			{9'd210, 8'd69}: color_data = 12'h09e;
			{9'd210, 8'd70}: color_data = 12'h09e;
			{9'd210, 8'd71}: color_data = 12'h09e;
			{9'd210, 8'd72}: color_data = 12'h09e;
			{9'd210, 8'd73}: color_data = 12'h09e;
			{9'd210, 8'd74}: color_data = 12'h09e;
			{9'd210, 8'd75}: color_data = 12'h09e;
			{9'd210, 8'd76}: color_data = 12'h08c;
			{9'd210, 8'd77}: color_data = 12'h023;
			{9'd210, 8'd119}: color_data = 12'h000;
			{9'd210, 8'd120}: color_data = 12'h07b;
			{9'd210, 8'd121}: color_data = 12'h0ae;
			{9'd210, 8'd122}: color_data = 12'h09e;
			{9'd210, 8'd123}: color_data = 12'h09e;
			{9'd210, 8'd124}: color_data = 12'h09e;
			{9'd210, 8'd125}: color_data = 12'h09e;
			{9'd210, 8'd126}: color_data = 12'h09e;
			{9'd210, 8'd127}: color_data = 12'h09e;
			{9'd210, 8'd128}: color_data = 12'h057;
			{9'd210, 8'd129}: color_data = 12'h000;
			{9'd210, 8'd170}: color_data = 12'h000;
			{9'd210, 8'd171}: color_data = 12'h057;
			{9'd210, 8'd172}: color_data = 12'h0ad;
			{9'd210, 8'd173}: color_data = 12'h09d;
			{9'd210, 8'd174}: color_data = 12'h09d;
			{9'd210, 8'd175}: color_data = 12'h09d;
			{9'd210, 8'd176}: color_data = 12'h09d;
			{9'd210, 8'd177}: color_data = 12'h09d;
			{9'd210, 8'd178}: color_data = 12'h09d;
			{9'd210, 8'd179}: color_data = 12'h08b;
			{9'd210, 8'd180}: color_data = 12'h012;
			{9'd210, 8'd222}: color_data = 12'h000;
			{9'd210, 8'd223}: color_data = 12'h200;
			{9'd210, 8'd224}: color_data = 12'h300;
			{9'd210, 8'd225}: color_data = 12'h100;
			{9'd210, 8'd226}: color_data = 12'h000;
			{9'd210, 8'd227}: color_data = 12'h700;
			{9'd210, 8'd228}: color_data = 12'ha00;
			{9'd210, 8'd229}: color_data = 12'h900;
			{9'd210, 8'd230}: color_data = 12'h300;
			{9'd210, 8'd231}: color_data = 12'h100;
			{9'd210, 8'd232}: color_data = 12'h310;
			{9'd210, 8'd233}: color_data = 12'h200;
			{9'd210, 8'd234}: color_data = 12'h000;
			{9'd210, 8'd235}: color_data = 12'h300;
			{9'd210, 8'd236}: color_data = 12'h900;
			{9'd210, 8'd237}: color_data = 12'ha00;
			{9'd210, 8'd238}: color_data = 12'h700;
			{9'd210, 8'd239}: color_data = 12'h100;
			{9'd211, 8'd68}: color_data = 12'h057;
			{9'd211, 8'd69}: color_data = 12'h4ef;
			{9'd211, 8'd70}: color_data = 12'h7ef;
			{9'd211, 8'd71}: color_data = 12'h0cf;
			{9'd211, 8'd72}: color_data = 12'h0cf;
			{9'd211, 8'd73}: color_data = 12'h0df;
			{9'd211, 8'd74}: color_data = 12'h0bd;
			{9'd211, 8'd75}: color_data = 12'h068;
			{9'd211, 8'd76}: color_data = 12'h09c;
			{9'd211, 8'd77}: color_data = 12'h034;
			{9'd211, 8'd119}: color_data = 12'h000;
			{9'd211, 8'd120}: color_data = 12'h1ad;
			{9'd211, 8'd121}: color_data = 12'h8ff;
			{9'd211, 8'd122}: color_data = 12'h3df;
			{9'd211, 8'd123}: color_data = 12'h0cf;
			{9'd211, 8'd124}: color_data = 12'h0cf;
			{9'd211, 8'd125}: color_data = 12'h0cf;
			{9'd211, 8'd126}: color_data = 12'h07a;
			{9'd211, 8'd127}: color_data = 12'h08b;
			{9'd211, 8'd128}: color_data = 12'h079;
			{9'd211, 8'd129}: color_data = 12'h000;
			{9'd211, 8'd170}: color_data = 12'h000;
			{9'd211, 8'd171}: color_data = 12'h069;
			{9'd211, 8'd172}: color_data = 12'h6ef;
			{9'd211, 8'd173}: color_data = 12'h6ef;
			{9'd211, 8'd174}: color_data = 12'h0cf;
			{9'd211, 8'd175}: color_data = 12'h0cf;
			{9'd211, 8'd176}: color_data = 12'h0df;
			{9'd211, 8'd177}: color_data = 12'h0ad;
			{9'd211, 8'd178}: color_data = 12'h079;
			{9'd211, 8'd179}: color_data = 12'h09c;
			{9'd211, 8'd180}: color_data = 12'h023;
			{9'd211, 8'd222}: color_data = 12'h100;
			{9'd211, 8'd223}: color_data = 12'h400;
			{9'd211, 8'd224}: color_data = 12'h500;
			{9'd211, 8'd225}: color_data = 12'h400;
			{9'd211, 8'd226}: color_data = 12'h200;
			{9'd211, 8'd227}: color_data = 12'ha20;
			{9'd211, 8'd228}: color_data = 12'hb10;
			{9'd211, 8'd229}: color_data = 12'h900;
			{9'd211, 8'd230}: color_data = 12'h300;
			{9'd211, 8'd231}: color_data = 12'h200;
			{9'd211, 8'd232}: color_data = 12'h500;
			{9'd211, 8'd233}: color_data = 12'h500;
			{9'd211, 8'd234}: color_data = 12'h200;
			{9'd211, 8'd235}: color_data = 12'h410;
			{9'd211, 8'd236}: color_data = 12'hc20;
			{9'd211, 8'd237}: color_data = 12'ha00;
			{9'd211, 8'd238}: color_data = 12'h700;
			{9'd211, 8'd239}: color_data = 12'h100;
			{9'd212, 8'd68}: color_data = 12'h047;
			{9'd212, 8'd69}: color_data = 12'h6df;
			{9'd212, 8'd70}: color_data = 12'heff;
			{9'd212, 8'd71}: color_data = 12'h6df;
			{9'd212, 8'd72}: color_data = 12'h0bf;
			{9'd212, 8'd73}: color_data = 12'h0be;
			{9'd212, 8'd74}: color_data = 12'h056;
			{9'd212, 8'd75}: color_data = 12'h012;
			{9'd212, 8'd76}: color_data = 12'h08b;
			{9'd212, 8'd77}: color_data = 12'h034;
			{9'd212, 8'd119}: color_data = 12'h000;
			{9'd212, 8'd120}: color_data = 12'h2ac;
			{9'd212, 8'd121}: color_data = 12'hdff;
			{9'd212, 8'd122}: color_data = 12'haef;
			{9'd212, 8'd123}: color_data = 12'h1cf;
			{9'd212, 8'd124}: color_data = 12'h0cf;
			{9'd212, 8'd125}: color_data = 12'h08b;
			{9'd212, 8'd126}: color_data = 12'h012;
			{9'd212, 8'd127}: color_data = 12'h068;
			{9'd212, 8'd128}: color_data = 12'h079;
			{9'd212, 8'd129}: color_data = 12'h000;
			{9'd212, 8'd170}: color_data = 12'h000;
			{9'd212, 8'd171}: color_data = 12'h068;
			{9'd212, 8'd172}: color_data = 12'h8ef;
			{9'd212, 8'd173}: color_data = 12'hdff;
			{9'd212, 8'd174}: color_data = 12'h4cf;
			{9'd212, 8'd175}: color_data = 12'h0bf;
			{9'd212, 8'd176}: color_data = 12'h0ae;
			{9'd212, 8'd177}: color_data = 12'h035;
			{9'd212, 8'd178}: color_data = 12'h023;
			{9'd212, 8'd179}: color_data = 12'h08c;
			{9'd212, 8'd180}: color_data = 12'h023;
			{9'd212, 8'd222}: color_data = 12'h200;
			{9'd212, 8'd223}: color_data = 12'h900;
			{9'd212, 8'd224}: color_data = 12'hb00;
			{9'd212, 8'd225}: color_data = 12'h800;
			{9'd212, 8'd226}: color_data = 12'h200;
			{9'd212, 8'd227}: color_data = 12'hb30;
			{9'd212, 8'd228}: color_data = 12'hc10;
			{9'd212, 8'd229}: color_data = 12'h800;
			{9'd212, 8'd230}: color_data = 12'h300;
			{9'd212, 8'd231}: color_data = 12'h400;
			{9'd212, 8'd232}: color_data = 12'ha00;
			{9'd212, 8'd233}: color_data = 12'ha00;
			{9'd212, 8'd234}: color_data = 12'h500;
			{9'd212, 8'd235}: color_data = 12'h510;
			{9'd212, 8'd236}: color_data = 12'hd30;
			{9'd212, 8'd237}: color_data = 12'ha00;
			{9'd212, 8'd238}: color_data = 12'h700;
			{9'd212, 8'd239}: color_data = 12'h100;
			{9'd213, 8'd68}: color_data = 12'h047;
			{9'd213, 8'd69}: color_data = 12'h6df;
			{9'd213, 8'd70}: color_data = 12'hfff;
			{9'd213, 8'd71}: color_data = 12'hdff;
			{9'd213, 8'd72}: color_data = 12'h5df;
			{9'd213, 8'd73}: color_data = 12'h068;
			{9'd213, 8'd74}: color_data = 12'h000;
			{9'd213, 8'd75}: color_data = 12'h012;
			{9'd213, 8'd76}: color_data = 12'h08c;
			{9'd213, 8'd77}: color_data = 12'h034;
			{9'd213, 8'd119}: color_data = 12'h000;
			{9'd213, 8'd120}: color_data = 12'h1ac;
			{9'd213, 8'd121}: color_data = 12'hdff;
			{9'd213, 8'd122}: color_data = 12'hfff;
			{9'd213, 8'd123}: color_data = 12'h9ef;
			{9'd213, 8'd124}: color_data = 12'h19c;
			{9'd213, 8'd125}: color_data = 12'h023;
			{9'd213, 8'd127}: color_data = 12'h068;
			{9'd213, 8'd128}: color_data = 12'h079;
			{9'd213, 8'd129}: color_data = 12'h000;
			{9'd213, 8'd170}: color_data = 12'h000;
			{9'd213, 8'd171}: color_data = 12'h068;
			{9'd213, 8'd172}: color_data = 12'h8ef;
			{9'd213, 8'd173}: color_data = 12'hfff;
			{9'd213, 8'd174}: color_data = 12'hcff;
			{9'd213, 8'd175}: color_data = 12'h4ce;
			{9'd213, 8'd176}: color_data = 12'h057;
			{9'd213, 8'd177}: color_data = 12'h000;
			{9'd213, 8'd178}: color_data = 12'h023;
			{9'd213, 8'd179}: color_data = 12'h08c;
			{9'd213, 8'd180}: color_data = 12'h023;
			{9'd213, 8'd222}: color_data = 12'h200;
			{9'd213, 8'd223}: color_data = 12'h900;
			{9'd213, 8'd224}: color_data = 12'ha00;
			{9'd213, 8'd225}: color_data = 12'h700;
			{9'd213, 8'd226}: color_data = 12'h200;
			{9'd213, 8'd227}: color_data = 12'hb30;
			{9'd213, 8'd228}: color_data = 12'he20;
			{9'd213, 8'd229}: color_data = 12'ha00;
			{9'd213, 8'd230}: color_data = 12'h300;
			{9'd213, 8'd231}: color_data = 12'h400;
			{9'd213, 8'd232}: color_data = 12'ha00;
			{9'd213, 8'd233}: color_data = 12'ha00;
			{9'd213, 8'd234}: color_data = 12'h400;
			{9'd213, 8'd235}: color_data = 12'h510;
			{9'd213, 8'd236}: color_data = 12'hf40;
			{9'd213, 8'd237}: color_data = 12'hd10;
			{9'd213, 8'd238}: color_data = 12'h800;
			{9'd213, 8'd239}: color_data = 12'h100;
			{9'd214, 8'd68}: color_data = 12'h047;
			{9'd214, 8'd69}: color_data = 12'h6df;
			{9'd214, 8'd70}: color_data = 12'hfff;
			{9'd214, 8'd71}: color_data = 12'hfff;
			{9'd214, 8'd72}: color_data = 12'h9aa;
			{9'd214, 8'd73}: color_data = 12'h011;
			{9'd214, 8'd75}: color_data = 12'h012;
			{9'd214, 8'd76}: color_data = 12'h08c;
			{9'd214, 8'd77}: color_data = 12'h034;
			{9'd214, 8'd119}: color_data = 12'h000;
			{9'd214, 8'd120}: color_data = 12'h1ac;
			{9'd214, 8'd121}: color_data = 12'hcff;
			{9'd214, 8'd122}: color_data = 12'hfff;
			{9'd214, 8'd123}: color_data = 12'hddd;
			{9'd214, 8'd124}: color_data = 12'h345;
			{9'd214, 8'd126}: color_data = 12'h000;
			{9'd214, 8'd127}: color_data = 12'h068;
			{9'd214, 8'd128}: color_data = 12'h079;
			{9'd214, 8'd129}: color_data = 12'h000;
			{9'd214, 8'd170}: color_data = 12'h000;
			{9'd214, 8'd171}: color_data = 12'h068;
			{9'd214, 8'd172}: color_data = 12'h7ef;
			{9'd214, 8'd173}: color_data = 12'hfff;
			{9'd214, 8'd174}: color_data = 12'hfff;
			{9'd214, 8'd175}: color_data = 12'h899;
			{9'd214, 8'd176}: color_data = 12'h001;
			{9'd214, 8'd178}: color_data = 12'h024;
			{9'd214, 8'd179}: color_data = 12'h08c;
			{9'd214, 8'd180}: color_data = 12'h023;
			{9'd214, 8'd222}: color_data = 12'h200;
			{9'd214, 8'd223}: color_data = 12'h800;
			{9'd214, 8'd224}: color_data = 12'ha00;
			{9'd214, 8'd225}: color_data = 12'h800;
			{9'd214, 8'd226}: color_data = 12'h200;
			{9'd214, 8'd227}: color_data = 12'h920;
			{9'd214, 8'd228}: color_data = 12'hd30;
			{9'd214, 8'd229}: color_data = 12'h910;
			{9'd214, 8'd230}: color_data = 12'h200;
			{9'd214, 8'd231}: color_data = 12'h400;
			{9'd214, 8'd232}: color_data = 12'h900;
			{9'd214, 8'd233}: color_data = 12'ha00;
			{9'd214, 8'd234}: color_data = 12'h400;
			{9'd214, 8'd235}: color_data = 12'h310;
			{9'd214, 8'd236}: color_data = 12'hc30;
			{9'd214, 8'd237}: color_data = 12'hc20;
			{9'd214, 8'd238}: color_data = 12'h600;
			{9'd214, 8'd239}: color_data = 12'h000;
			{9'd215, 8'd68}: color_data = 12'h047;
			{9'd215, 8'd69}: color_data = 12'h6df;
			{9'd215, 8'd70}: color_data = 12'hfff;
			{9'd215, 8'd71}: color_data = 12'hcbb;
			{9'd215, 8'd72}: color_data = 12'h323;
			{9'd215, 8'd73}: color_data = 12'h002;
			{9'd215, 8'd74}: color_data = 12'h000;
			{9'd215, 8'd75}: color_data = 12'h012;
			{9'd215, 8'd76}: color_data = 12'h08c;
			{9'd215, 8'd77}: color_data = 12'h034;
			{9'd215, 8'd119}: color_data = 12'h000;
			{9'd215, 8'd120}: color_data = 12'h1ac;
			{9'd215, 8'd121}: color_data = 12'hdff;
			{9'd215, 8'd122}: color_data = 12'hfee;
			{9'd215, 8'd123}: color_data = 12'h666;
			{9'd215, 8'd124}: color_data = 12'h002;
			{9'd215, 8'd125}: color_data = 12'h001;
			{9'd215, 8'd126}: color_data = 12'h000;
			{9'd215, 8'd127}: color_data = 12'h068;
			{9'd215, 8'd128}: color_data = 12'h079;
			{9'd215, 8'd129}: color_data = 12'h000;
			{9'd215, 8'd170}: color_data = 12'h000;
			{9'd215, 8'd171}: color_data = 12'h068;
			{9'd215, 8'd172}: color_data = 12'h8ef;
			{9'd215, 8'd173}: color_data = 12'hfff;
			{9'd215, 8'd174}: color_data = 12'haa9;
			{9'd215, 8'd175}: color_data = 12'h212;
			{9'd215, 8'd176}: color_data = 12'h002;
			{9'd215, 8'd177}: color_data = 12'h000;
			{9'd215, 8'd178}: color_data = 12'h023;
			{9'd215, 8'd179}: color_data = 12'h08c;
			{9'd215, 8'd180}: color_data = 12'h023;
			{9'd215, 8'd222}: color_data = 12'h200;
			{9'd215, 8'd223}: color_data = 12'h900;
			{9'd215, 8'd224}: color_data = 12'ha00;
			{9'd215, 8'd225}: color_data = 12'h800;
			{9'd215, 8'd226}: color_data = 12'h100;
			{9'd215, 8'd227}: color_data = 12'h100;
			{9'd215, 8'd228}: color_data = 12'h310;
			{9'd215, 8'd229}: color_data = 12'h200;
			{9'd215, 8'd230}: color_data = 12'h000;
			{9'd215, 8'd231}: color_data = 12'h500;
			{9'd215, 8'd232}: color_data = 12'ha00;
			{9'd215, 8'd233}: color_data = 12'ha00;
			{9'd215, 8'd234}: color_data = 12'h500;
			{9'd215, 8'd235}: color_data = 12'h000;
			{9'd215, 8'd236}: color_data = 12'h200;
			{9'd215, 8'd237}: color_data = 12'h300;
			{9'd215, 8'd238}: color_data = 12'h100;
			{9'd215, 8'd239}: color_data = 12'h000;
			{9'd216, 8'd68}: color_data = 12'h047;
			{9'd216, 8'd69}: color_data = 12'h6ef;
			{9'd216, 8'd70}: color_data = 12'hccc;
			{9'd216, 8'd71}: color_data = 12'h434;
			{9'd216, 8'd72}: color_data = 12'h003;
			{9'd216, 8'd73}: color_data = 12'h005;
			{9'd216, 8'd74}: color_data = 12'h002;
			{9'd216, 8'd75}: color_data = 12'h012;
			{9'd216, 8'd76}: color_data = 12'h08c;
			{9'd216, 8'd77}: color_data = 12'h034;
			{9'd216, 8'd119}: color_data = 12'h000;
			{9'd216, 8'd120}: color_data = 12'h2ad;
			{9'd216, 8'd121}: color_data = 12'hcff;
			{9'd216, 8'd122}: color_data = 12'h877;
			{9'd216, 8'd123}: color_data = 12'h002;
			{9'd216, 8'd124}: color_data = 12'h004;
			{9'd216, 8'd125}: color_data = 12'h004;
			{9'd216, 8'd126}: color_data = 12'h000;
			{9'd216, 8'd127}: color_data = 12'h068;
			{9'd216, 8'd128}: color_data = 12'h079;
			{9'd216, 8'd129}: color_data = 12'h000;
			{9'd216, 8'd170}: color_data = 12'h000;
			{9'd216, 8'd171}: color_data = 12'h068;
			{9'd216, 8'd172}: color_data = 12'h8ff;
			{9'd216, 8'd173}: color_data = 12'hcbb;
			{9'd216, 8'd174}: color_data = 12'h223;
			{9'd216, 8'd175}: color_data = 12'h003;
			{9'd216, 8'd176}: color_data = 12'h005;
			{9'd216, 8'd177}: color_data = 12'h002;
			{9'd216, 8'd178}: color_data = 12'h023;
			{9'd216, 8'd179}: color_data = 12'h09c;
			{9'd216, 8'd180}: color_data = 12'h023;
			{9'd216, 8'd222}: color_data = 12'h300;
			{9'd216, 8'd223}: color_data = 12'hc20;
			{9'd216, 8'd224}: color_data = 12'ha00;
			{9'd216, 8'd225}: color_data = 12'h800;
			{9'd216, 8'd226}: color_data = 12'h100;
			{9'd216, 8'd227}: color_data = 12'h300;
			{9'd216, 8'd228}: color_data = 12'h500;
			{9'd216, 8'd229}: color_data = 12'h500;
			{9'd216, 8'd230}: color_data = 12'h100;
			{9'd216, 8'd231}: color_data = 12'h710;
			{9'd216, 8'd232}: color_data = 12'hc10;
			{9'd216, 8'd233}: color_data = 12'h900;
			{9'd216, 8'd234}: color_data = 12'h500;
			{9'd216, 8'd235}: color_data = 12'h100;
			{9'd216, 8'd236}: color_data = 12'h500;
			{9'd216, 8'd237}: color_data = 12'h500;
			{9'd216, 8'd238}: color_data = 12'h400;
			{9'd216, 8'd239}: color_data = 12'h000;
			{9'd217, 8'd68}: color_data = 12'h057;
			{9'd217, 8'd69}: color_data = 12'h3bd;
			{9'd217, 8'd70}: color_data = 12'h555;
			{9'd217, 8'd71}: color_data = 12'h002;
			{9'd217, 8'd72}: color_data = 12'h005;
			{9'd217, 8'd73}: color_data = 12'h005;
			{9'd217, 8'd74}: color_data = 12'h004;
			{9'd217, 8'd75}: color_data = 12'h025;
			{9'd217, 8'd76}: color_data = 12'h09c;
			{9'd217, 8'd77}: color_data = 12'h034;
			{9'd217, 8'd119}: color_data = 12'h000;
			{9'd217, 8'd120}: color_data = 12'h1ac;
			{9'd217, 8'd121}: color_data = 12'h689;
			{9'd217, 8'd122}: color_data = 12'h212;
			{9'd217, 8'd123}: color_data = 12'h004;
			{9'd217, 8'd124}: color_data = 12'h005;
			{9'd217, 8'd125}: color_data = 12'h005;
			{9'd217, 8'd126}: color_data = 12'h003;
			{9'd217, 8'd127}: color_data = 12'h06a;
			{9'd217, 8'd128}: color_data = 12'h079;
			{9'd217, 8'd129}: color_data = 12'h000;
			{9'd217, 8'd170}: color_data = 12'h000;
			{9'd217, 8'd171}: color_data = 12'h079;
			{9'd217, 8'd172}: color_data = 12'h4bd;
			{9'd217, 8'd173}: color_data = 12'h444;
			{9'd217, 8'd174}: color_data = 12'h002;
			{9'd217, 8'd175}: color_data = 12'h005;
			{9'd217, 8'd176}: color_data = 12'h005;
			{9'd217, 8'd177}: color_data = 12'h004;
			{9'd217, 8'd178}: color_data = 12'h036;
			{9'd217, 8'd179}: color_data = 12'h09c;
			{9'd217, 8'd180}: color_data = 12'h023;
			{9'd217, 8'd222}: color_data = 12'h410;
			{9'd217, 8'd223}: color_data = 12'hd30;
			{9'd217, 8'd224}: color_data = 12'hb00;
			{9'd217, 8'd225}: color_data = 12'h700;
			{9'd217, 8'd226}: color_data = 12'h200;
			{9'd217, 8'd227}: color_data = 12'h700;
			{9'd217, 8'd228}: color_data = 12'hb00;
			{9'd217, 8'd229}: color_data = 12'ha00;
			{9'd217, 8'd230}: color_data = 12'h300;
			{9'd217, 8'd231}: color_data = 12'h820;
			{9'd217, 8'd232}: color_data = 12'hd20;
			{9'd217, 8'd233}: color_data = 12'h900;
			{9'd217, 8'd234}: color_data = 12'h500;
			{9'd217, 8'd235}: color_data = 12'h300;
			{9'd217, 8'd236}: color_data = 12'h900;
			{9'd217, 8'd237}: color_data = 12'hb00;
			{9'd217, 8'd238}: color_data = 12'h800;
			{9'd217, 8'd239}: color_data = 12'h100;
			{9'd218, 8'd68}: color_data = 12'h035;
			{9'd218, 8'd69}: color_data = 12'h047;
			{9'd218, 8'd70}: color_data = 12'h001;
			{9'd218, 8'd71}: color_data = 12'h004;
			{9'd218, 8'd72}: color_data = 12'h004;
			{9'd218, 8'd73}: color_data = 12'h004;
			{9'd218, 8'd74}: color_data = 12'h004;
			{9'd218, 8'd75}: color_data = 12'h015;
			{9'd218, 8'd76}: color_data = 12'h059;
			{9'd218, 8'd77}: color_data = 12'h023;
			{9'd218, 8'd119}: color_data = 12'h000;
			{9'd218, 8'd120}: color_data = 12'h058;
			{9'd218, 8'd121}: color_data = 12'h013;
			{9'd218, 8'd122}: color_data = 12'h002;
			{9'd218, 8'd123}: color_data = 12'h004;
			{9'd218, 8'd124}: color_data = 12'h004;
			{9'd218, 8'd125}: color_data = 12'h004;
			{9'd218, 8'd126}: color_data = 12'h004;
			{9'd218, 8'd127}: color_data = 12'h038;
			{9'd218, 8'd128}: color_data = 12'h046;
			{9'd218, 8'd129}: color_data = 12'h000;
			{9'd218, 8'd170}: color_data = 12'h000;
			{9'd218, 8'd171}: color_data = 12'h047;
			{9'd218, 8'd172}: color_data = 12'h036;
			{9'd218, 8'd173}: color_data = 12'h001;
			{9'd218, 8'd174}: color_data = 12'h004;
			{9'd218, 8'd175}: color_data = 12'h004;
			{9'd218, 8'd176}: color_data = 12'h004;
			{9'd218, 8'd177}: color_data = 12'h004;
			{9'd218, 8'd178}: color_data = 12'h016;
			{9'd218, 8'd179}: color_data = 12'h059;
			{9'd218, 8'd180}: color_data = 12'h012;
			{9'd218, 8'd222}: color_data = 12'h410;
			{9'd218, 8'd223}: color_data = 12'he40;
			{9'd218, 8'd224}: color_data = 12'hd20;
			{9'd218, 8'd225}: color_data = 12'h800;
			{9'd218, 8'd226}: color_data = 12'h200;
			{9'd218, 8'd227}: color_data = 12'h600;
			{9'd218, 8'd228}: color_data = 12'ha00;
			{9'd218, 8'd229}: color_data = 12'h900;
			{9'd218, 8'd230}: color_data = 12'h300;
			{9'd218, 8'd231}: color_data = 12'h820;
			{9'd218, 8'd232}: color_data = 12'hf30;
			{9'd218, 8'd233}: color_data = 12'hc00;
			{9'd218, 8'd234}: color_data = 12'h500;
			{9'd218, 8'd235}: color_data = 12'h200;
			{9'd218, 8'd236}: color_data = 12'h900;
			{9'd218, 8'd237}: color_data = 12'ha00;
			{9'd218, 8'd238}: color_data = 12'h700;
			{9'd218, 8'd239}: color_data = 12'h100;
			{9'd219, 8'd68}: color_data = 12'h013;
			{9'd219, 8'd69}: color_data = 12'h027;
			{9'd219, 8'd70}: color_data = 12'h016;
			{9'd219, 8'd71}: color_data = 12'h027;
			{9'd219, 8'd72}: color_data = 12'h027;
			{9'd219, 8'd73}: color_data = 12'h027;
			{9'd219, 8'd74}: color_data = 12'h027;
			{9'd219, 8'd75}: color_data = 12'h028;
			{9'd219, 8'd76}: color_data = 12'h027;
			{9'd219, 8'd77}: color_data = 12'h001;
			{9'd219, 8'd119}: color_data = 12'h000;
			{9'd219, 8'd120}: color_data = 12'h016;
			{9'd219, 8'd121}: color_data = 12'h017;
			{9'd219, 8'd122}: color_data = 12'h016;
			{9'd219, 8'd123}: color_data = 12'h027;
			{9'd219, 8'd124}: color_data = 12'h027;
			{9'd219, 8'd125}: color_data = 12'h027;
			{9'd219, 8'd126}: color_data = 12'h027;
			{9'd219, 8'd127}: color_data = 12'h028;
			{9'd219, 8'd128}: color_data = 12'h014;
			{9'd219, 8'd129}: color_data = 12'h000;
			{9'd219, 8'd170}: color_data = 12'h000;
			{9'd219, 8'd171}: color_data = 12'h014;
			{9'd219, 8'd172}: color_data = 12'h027;
			{9'd219, 8'd173}: color_data = 12'h016;
			{9'd219, 8'd174}: color_data = 12'h027;
			{9'd219, 8'd175}: color_data = 12'h027;
			{9'd219, 8'd176}: color_data = 12'h027;
			{9'd219, 8'd177}: color_data = 12'h027;
			{9'd219, 8'd178}: color_data = 12'h028;
			{9'd219, 8'd179}: color_data = 12'h026;
			{9'd219, 8'd180}: color_data = 12'h001;
			{9'd219, 8'd222}: color_data = 12'h300;
			{9'd219, 8'd223}: color_data = 12'hc30;
			{9'd219, 8'd224}: color_data = 12'hc30;
			{9'd219, 8'd225}: color_data = 12'h700;
			{9'd219, 8'd226}: color_data = 12'h100;
			{9'd219, 8'd227}: color_data = 12'h600;
			{9'd219, 8'd228}: color_data = 12'ha00;
			{9'd219, 8'd229}: color_data = 12'h900;
			{9'd219, 8'd230}: color_data = 12'h300;
			{9'd219, 8'd231}: color_data = 12'h620;
			{9'd219, 8'd232}: color_data = 12'hd40;
			{9'd219, 8'd233}: color_data = 12'ha20;
			{9'd219, 8'd234}: color_data = 12'h300;
			{9'd219, 8'd235}: color_data = 12'h200;
			{9'd219, 8'd236}: color_data = 12'h900;
			{9'd219, 8'd237}: color_data = 12'ha00;
			{9'd219, 8'd238}: color_data = 12'h700;
			{9'd219, 8'd239}: color_data = 12'h100;
			{9'd220, 8'd68}: color_data = 12'h035;
			{9'd220, 8'd69}: color_data = 12'h09e;
			{9'd220, 8'd70}: color_data = 12'h09e;
			{9'd220, 8'd71}: color_data = 12'h09e;
			{9'd220, 8'd72}: color_data = 12'h09e;
			{9'd220, 8'd73}: color_data = 12'h09e;
			{9'd220, 8'd74}: color_data = 12'h09e;
			{9'd220, 8'd75}: color_data = 12'h09e;
			{9'd220, 8'd76}: color_data = 12'h08c;
			{9'd220, 8'd77}: color_data = 12'h023;
			{9'd220, 8'd119}: color_data = 12'h000;
			{9'd220, 8'd120}: color_data = 12'h07b;
			{9'd220, 8'd121}: color_data = 12'h0ae;
			{9'd220, 8'd122}: color_data = 12'h09e;
			{9'd220, 8'd123}: color_data = 12'h09e;
			{9'd220, 8'd124}: color_data = 12'h09e;
			{9'd220, 8'd125}: color_data = 12'h09e;
			{9'd220, 8'd126}: color_data = 12'h09e;
			{9'd220, 8'd127}: color_data = 12'h09e;
			{9'd220, 8'd128}: color_data = 12'h057;
			{9'd220, 8'd129}: color_data = 12'h000;
			{9'd220, 8'd170}: color_data = 12'h000;
			{9'd220, 8'd171}: color_data = 12'h057;
			{9'd220, 8'd172}: color_data = 12'h0ae;
			{9'd220, 8'd173}: color_data = 12'h09e;
			{9'd220, 8'd174}: color_data = 12'h09e;
			{9'd220, 8'd175}: color_data = 12'h09e;
			{9'd220, 8'd176}: color_data = 12'h09e;
			{9'd220, 8'd177}: color_data = 12'h09e;
			{9'd220, 8'd178}: color_data = 12'h09e;
			{9'd220, 8'd179}: color_data = 12'h07b;
			{9'd220, 8'd180}: color_data = 12'h012;
			{9'd220, 8'd222}: color_data = 12'h000;
			{9'd220, 8'd223}: color_data = 12'h200;
			{9'd220, 8'd224}: color_data = 12'h300;
			{9'd220, 8'd225}: color_data = 12'h100;
			{9'd220, 8'd226}: color_data = 12'h000;
			{9'd220, 8'd227}: color_data = 12'h700;
			{9'd220, 8'd228}: color_data = 12'ha00;
			{9'd220, 8'd229}: color_data = 12'h900;
			{9'd220, 8'd230}: color_data = 12'h300;
			{9'd220, 8'd231}: color_data = 12'h100;
			{9'd220, 8'd232}: color_data = 12'h310;
			{9'd220, 8'd233}: color_data = 12'h200;
			{9'd220, 8'd234}: color_data = 12'h000;
			{9'd220, 8'd235}: color_data = 12'h300;
			{9'd220, 8'd236}: color_data = 12'h900;
			{9'd220, 8'd237}: color_data = 12'ha00;
			{9'd220, 8'd238}: color_data = 12'h700;
			{9'd220, 8'd239}: color_data = 12'h100;
			{9'd221, 8'd68}: color_data = 12'h057;
			{9'd221, 8'd69}: color_data = 12'h4ef;
			{9'd221, 8'd70}: color_data = 12'h7ef;
			{9'd221, 8'd71}: color_data = 12'h0cf;
			{9'd221, 8'd72}: color_data = 12'h0cf;
			{9'd221, 8'd73}: color_data = 12'h0df;
			{9'd221, 8'd74}: color_data = 12'h0bd;
			{9'd221, 8'd75}: color_data = 12'h068;
			{9'd221, 8'd76}: color_data = 12'h09c;
			{9'd221, 8'd77}: color_data = 12'h034;
			{9'd221, 8'd119}: color_data = 12'h000;
			{9'd221, 8'd120}: color_data = 12'h1ad;
			{9'd221, 8'd121}: color_data = 12'h8ff;
			{9'd221, 8'd122}: color_data = 12'h3df;
			{9'd221, 8'd123}: color_data = 12'h0bf;
			{9'd221, 8'd124}: color_data = 12'h0cf;
			{9'd221, 8'd125}: color_data = 12'h0cf;
			{9'd221, 8'd126}: color_data = 12'h079;
			{9'd221, 8'd127}: color_data = 12'h08b;
			{9'd221, 8'd128}: color_data = 12'h079;
			{9'd221, 8'd129}: color_data = 12'h000;
			{9'd221, 8'd170}: color_data = 12'h000;
			{9'd221, 8'd171}: color_data = 12'h069;
			{9'd221, 8'd172}: color_data = 12'h6ef;
			{9'd221, 8'd173}: color_data = 12'h6ef;
			{9'd221, 8'd174}: color_data = 12'h0cf;
			{9'd221, 8'd175}: color_data = 12'h0cf;
			{9'd221, 8'd176}: color_data = 12'h0df;
			{9'd221, 8'd177}: color_data = 12'h0ac;
			{9'd221, 8'd178}: color_data = 12'h079;
			{9'd221, 8'd179}: color_data = 12'h09c;
			{9'd221, 8'd180}: color_data = 12'h023;
			{9'd221, 8'd222}: color_data = 12'h100;
			{9'd221, 8'd223}: color_data = 12'h500;
			{9'd221, 8'd224}: color_data = 12'h500;
			{9'd221, 8'd225}: color_data = 12'h400;
			{9'd221, 8'd226}: color_data = 12'h200;
			{9'd221, 8'd227}: color_data = 12'ha20;
			{9'd221, 8'd228}: color_data = 12'hb10;
			{9'd221, 8'd229}: color_data = 12'h900;
			{9'd221, 8'd230}: color_data = 12'h300;
			{9'd221, 8'd231}: color_data = 12'h200;
			{9'd221, 8'd232}: color_data = 12'h500;
			{9'd221, 8'd233}: color_data = 12'h500;
			{9'd221, 8'd234}: color_data = 12'h200;
			{9'd221, 8'd235}: color_data = 12'h410;
			{9'd221, 8'd236}: color_data = 12'hc20;
			{9'd221, 8'd237}: color_data = 12'ha00;
			{9'd221, 8'd238}: color_data = 12'h700;
			{9'd221, 8'd239}: color_data = 12'h100;
			{9'd222, 8'd68}: color_data = 12'h047;
			{9'd222, 8'd69}: color_data = 12'h6df;
			{9'd222, 8'd70}: color_data = 12'heff;
			{9'd222, 8'd71}: color_data = 12'h6df;
			{9'd222, 8'd72}: color_data = 12'h0bf;
			{9'd222, 8'd73}: color_data = 12'h0bf;
			{9'd222, 8'd74}: color_data = 12'h056;
			{9'd222, 8'd75}: color_data = 12'h012;
			{9'd222, 8'd76}: color_data = 12'h08b;
			{9'd222, 8'd77}: color_data = 12'h034;
			{9'd222, 8'd119}: color_data = 12'h000;
			{9'd222, 8'd120}: color_data = 12'h2ac;
			{9'd222, 8'd121}: color_data = 12'hdff;
			{9'd222, 8'd122}: color_data = 12'haef;
			{9'd222, 8'd123}: color_data = 12'h1bf;
			{9'd222, 8'd124}: color_data = 12'h0cf;
			{9'd222, 8'd125}: color_data = 12'h08b;
			{9'd222, 8'd126}: color_data = 12'h012;
			{9'd222, 8'd127}: color_data = 12'h058;
			{9'd222, 8'd128}: color_data = 12'h079;
			{9'd222, 8'd129}: color_data = 12'h000;
			{9'd222, 8'd170}: color_data = 12'h000;
			{9'd222, 8'd171}: color_data = 12'h068;
			{9'd222, 8'd172}: color_data = 12'h8ef;
			{9'd222, 8'd173}: color_data = 12'hdff;
			{9'd222, 8'd174}: color_data = 12'h4cf;
			{9'd222, 8'd175}: color_data = 12'h0bf;
			{9'd222, 8'd176}: color_data = 12'h0ae;
			{9'd222, 8'd177}: color_data = 12'h035;
			{9'd222, 8'd178}: color_data = 12'h023;
			{9'd222, 8'd179}: color_data = 12'h08c;
			{9'd222, 8'd180}: color_data = 12'h023;
			{9'd222, 8'd222}: color_data = 12'h200;
			{9'd222, 8'd223}: color_data = 12'h900;
			{9'd222, 8'd224}: color_data = 12'hb00;
			{9'd222, 8'd225}: color_data = 12'h800;
			{9'd222, 8'd226}: color_data = 12'h200;
			{9'd222, 8'd227}: color_data = 12'hb30;
			{9'd222, 8'd228}: color_data = 12'hc10;
			{9'd222, 8'd229}: color_data = 12'h800;
			{9'd222, 8'd230}: color_data = 12'h300;
			{9'd222, 8'd231}: color_data = 12'h400;
			{9'd222, 8'd232}: color_data = 12'ha00;
			{9'd222, 8'd233}: color_data = 12'ha00;
			{9'd222, 8'd234}: color_data = 12'h500;
			{9'd222, 8'd235}: color_data = 12'h510;
			{9'd222, 8'd236}: color_data = 12'hd30;
			{9'd222, 8'd237}: color_data = 12'ha00;
			{9'd222, 8'd238}: color_data = 12'h700;
			{9'd222, 8'd239}: color_data = 12'h100;
			{9'd223, 8'd68}: color_data = 12'h047;
			{9'd223, 8'd69}: color_data = 12'h6df;
			{9'd223, 8'd70}: color_data = 12'hfff;
			{9'd223, 8'd71}: color_data = 12'hdff;
			{9'd223, 8'd72}: color_data = 12'h5df;
			{9'd223, 8'd73}: color_data = 12'h068;
			{9'd223, 8'd74}: color_data = 12'h000;
			{9'd223, 8'd75}: color_data = 12'h012;
			{9'd223, 8'd76}: color_data = 12'h08c;
			{9'd223, 8'd77}: color_data = 12'h034;
			{9'd223, 8'd119}: color_data = 12'h000;
			{9'd223, 8'd120}: color_data = 12'h1ac;
			{9'd223, 8'd121}: color_data = 12'hdff;
			{9'd223, 8'd122}: color_data = 12'hfff;
			{9'd223, 8'd123}: color_data = 12'h9ef;
			{9'd223, 8'd124}: color_data = 12'h19c;
			{9'd223, 8'd125}: color_data = 12'h023;
			{9'd223, 8'd127}: color_data = 12'h068;
			{9'd223, 8'd128}: color_data = 12'h079;
			{9'd223, 8'd129}: color_data = 12'h000;
			{9'd223, 8'd170}: color_data = 12'h000;
			{9'd223, 8'd171}: color_data = 12'h068;
			{9'd223, 8'd172}: color_data = 12'h8ef;
			{9'd223, 8'd173}: color_data = 12'hfff;
			{9'd223, 8'd174}: color_data = 12'hcff;
			{9'd223, 8'd175}: color_data = 12'h4ce;
			{9'd223, 8'd176}: color_data = 12'h057;
			{9'd223, 8'd177}: color_data = 12'h000;
			{9'd223, 8'd178}: color_data = 12'h023;
			{9'd223, 8'd179}: color_data = 12'h08c;
			{9'd223, 8'd180}: color_data = 12'h023;
			{9'd223, 8'd222}: color_data = 12'h200;
			{9'd223, 8'd223}: color_data = 12'h900;
			{9'd223, 8'd224}: color_data = 12'ha00;
			{9'd223, 8'd225}: color_data = 12'h700;
			{9'd223, 8'd226}: color_data = 12'h200;
			{9'd223, 8'd227}: color_data = 12'hb30;
			{9'd223, 8'd228}: color_data = 12'he20;
			{9'd223, 8'd229}: color_data = 12'ha00;
			{9'd223, 8'd230}: color_data = 12'h300;
			{9'd223, 8'd231}: color_data = 12'h400;
			{9'd223, 8'd232}: color_data = 12'ha00;
			{9'd223, 8'd233}: color_data = 12'ha00;
			{9'd223, 8'd234}: color_data = 12'h400;
			{9'd223, 8'd235}: color_data = 12'h510;
			{9'd223, 8'd236}: color_data = 12'hf40;
			{9'd223, 8'd237}: color_data = 12'hd10;
			{9'd223, 8'd238}: color_data = 12'h800;
			{9'd223, 8'd239}: color_data = 12'h100;
			{9'd224, 8'd68}: color_data = 12'h047;
			{9'd224, 8'd69}: color_data = 12'h6df;
			{9'd224, 8'd70}: color_data = 12'hfff;
			{9'd224, 8'd71}: color_data = 12'hfff;
			{9'd224, 8'd72}: color_data = 12'h9aa;
			{9'd224, 8'd73}: color_data = 12'h011;
			{9'd224, 8'd75}: color_data = 12'h012;
			{9'd224, 8'd76}: color_data = 12'h08c;
			{9'd224, 8'd77}: color_data = 12'h034;
			{9'd224, 8'd119}: color_data = 12'h000;
			{9'd224, 8'd120}: color_data = 12'h1ac;
			{9'd224, 8'd121}: color_data = 12'hcff;
			{9'd224, 8'd122}: color_data = 12'hfff;
			{9'd224, 8'd123}: color_data = 12'hddd;
			{9'd224, 8'd124}: color_data = 12'h345;
			{9'd224, 8'd126}: color_data = 12'h000;
			{9'd224, 8'd127}: color_data = 12'h068;
			{9'd224, 8'd128}: color_data = 12'h079;
			{9'd224, 8'd129}: color_data = 12'h000;
			{9'd224, 8'd170}: color_data = 12'h000;
			{9'd224, 8'd171}: color_data = 12'h068;
			{9'd224, 8'd172}: color_data = 12'h7ef;
			{9'd224, 8'd173}: color_data = 12'hfff;
			{9'd224, 8'd174}: color_data = 12'hfff;
			{9'd224, 8'd175}: color_data = 12'h899;
			{9'd224, 8'd176}: color_data = 12'h001;
			{9'd224, 8'd178}: color_data = 12'h024;
			{9'd224, 8'd179}: color_data = 12'h08c;
			{9'd224, 8'd180}: color_data = 12'h023;
			{9'd224, 8'd222}: color_data = 12'h200;
			{9'd224, 8'd223}: color_data = 12'h800;
			{9'd224, 8'd224}: color_data = 12'ha00;
			{9'd224, 8'd225}: color_data = 12'h700;
			{9'd224, 8'd226}: color_data = 12'h200;
			{9'd224, 8'd227}: color_data = 12'h920;
			{9'd224, 8'd228}: color_data = 12'hd30;
			{9'd224, 8'd229}: color_data = 12'h910;
			{9'd224, 8'd230}: color_data = 12'h200;
			{9'd224, 8'd231}: color_data = 12'h400;
			{9'd224, 8'd232}: color_data = 12'h900;
			{9'd224, 8'd233}: color_data = 12'ha00;
			{9'd224, 8'd234}: color_data = 12'h400;
			{9'd224, 8'd235}: color_data = 12'h310;
			{9'd224, 8'd236}: color_data = 12'hc30;
			{9'd224, 8'd237}: color_data = 12'hc20;
			{9'd224, 8'd238}: color_data = 12'h600;
			{9'd224, 8'd239}: color_data = 12'h000;
			{9'd225, 8'd68}: color_data = 12'h047;
			{9'd225, 8'd69}: color_data = 12'h6df;
			{9'd225, 8'd70}: color_data = 12'hfff;
			{9'd225, 8'd71}: color_data = 12'hcbb;
			{9'd225, 8'd72}: color_data = 12'h323;
			{9'd225, 8'd73}: color_data = 12'h002;
			{9'd225, 8'd74}: color_data = 12'h000;
			{9'd225, 8'd75}: color_data = 12'h012;
			{9'd225, 8'd76}: color_data = 12'h08c;
			{9'd225, 8'd77}: color_data = 12'h034;
			{9'd225, 8'd119}: color_data = 12'h000;
			{9'd225, 8'd120}: color_data = 12'h1ac;
			{9'd225, 8'd121}: color_data = 12'hdff;
			{9'd225, 8'd122}: color_data = 12'hfee;
			{9'd225, 8'd123}: color_data = 12'h666;
			{9'd225, 8'd124}: color_data = 12'h002;
			{9'd225, 8'd125}: color_data = 12'h001;
			{9'd225, 8'd126}: color_data = 12'h000;
			{9'd225, 8'd127}: color_data = 12'h068;
			{9'd225, 8'd128}: color_data = 12'h079;
			{9'd225, 8'd129}: color_data = 12'h000;
			{9'd225, 8'd170}: color_data = 12'h000;
			{9'd225, 8'd171}: color_data = 12'h068;
			{9'd225, 8'd172}: color_data = 12'h8ef;
			{9'd225, 8'd173}: color_data = 12'hfff;
			{9'd225, 8'd174}: color_data = 12'haaa;
			{9'd225, 8'd175}: color_data = 12'h213;
			{9'd225, 8'd176}: color_data = 12'h002;
			{9'd225, 8'd178}: color_data = 12'h023;
			{9'd225, 8'd179}: color_data = 12'h08c;
			{9'd225, 8'd180}: color_data = 12'h023;
			{9'd225, 8'd222}: color_data = 12'h200;
			{9'd225, 8'd223}: color_data = 12'h900;
			{9'd225, 8'd224}: color_data = 12'ha00;
			{9'd225, 8'd225}: color_data = 12'h800;
			{9'd225, 8'd226}: color_data = 12'h100;
			{9'd225, 8'd227}: color_data = 12'h100;
			{9'd225, 8'd228}: color_data = 12'h310;
			{9'd225, 8'd229}: color_data = 12'h200;
			{9'd225, 8'd230}: color_data = 12'h000;
			{9'd225, 8'd231}: color_data = 12'h500;
			{9'd225, 8'd232}: color_data = 12'ha00;
			{9'd225, 8'd233}: color_data = 12'ha00;
			{9'd225, 8'd234}: color_data = 12'h500;
			{9'd225, 8'd235}: color_data = 12'h000;
			{9'd225, 8'd236}: color_data = 12'h200;
			{9'd225, 8'd237}: color_data = 12'h300;
			{9'd225, 8'd238}: color_data = 12'h100;
			{9'd225, 8'd239}: color_data = 12'h000;
			{9'd226, 8'd68}: color_data = 12'h047;
			{9'd226, 8'd69}: color_data = 12'h6ef;
			{9'd226, 8'd70}: color_data = 12'hddc;
			{9'd226, 8'd71}: color_data = 12'h434;
			{9'd226, 8'd72}: color_data = 12'h003;
			{9'd226, 8'd73}: color_data = 12'h005;
			{9'd226, 8'd74}: color_data = 12'h002;
			{9'd226, 8'd75}: color_data = 12'h012;
			{9'd226, 8'd76}: color_data = 12'h08c;
			{9'd226, 8'd77}: color_data = 12'h034;
			{9'd226, 8'd119}: color_data = 12'h000;
			{9'd226, 8'd120}: color_data = 12'h2ad;
			{9'd226, 8'd121}: color_data = 12'hcff;
			{9'd226, 8'd122}: color_data = 12'h877;
			{9'd226, 8'd123}: color_data = 12'h002;
			{9'd226, 8'd124}: color_data = 12'h004;
			{9'd226, 8'd125}: color_data = 12'h004;
			{9'd226, 8'd126}: color_data = 12'h000;
			{9'd226, 8'd127}: color_data = 12'h068;
			{9'd226, 8'd128}: color_data = 12'h079;
			{9'd226, 8'd129}: color_data = 12'h000;
			{9'd226, 8'd170}: color_data = 12'h000;
			{9'd226, 8'd171}: color_data = 12'h068;
			{9'd226, 8'd172}: color_data = 12'h8ff;
			{9'd226, 8'd173}: color_data = 12'hcbb;
			{9'd226, 8'd174}: color_data = 12'h223;
			{9'd226, 8'd175}: color_data = 12'h003;
			{9'd226, 8'd176}: color_data = 12'h005;
			{9'd226, 8'd177}: color_data = 12'h002;
			{9'd226, 8'd178}: color_data = 12'h023;
			{9'd226, 8'd179}: color_data = 12'h09c;
			{9'd226, 8'd180}: color_data = 12'h023;
			{9'd226, 8'd222}: color_data = 12'h300;
			{9'd226, 8'd223}: color_data = 12'hc20;
			{9'd226, 8'd224}: color_data = 12'ha00;
			{9'd226, 8'd225}: color_data = 12'h800;
			{9'd226, 8'd226}: color_data = 12'h100;
			{9'd226, 8'd227}: color_data = 12'h300;
			{9'd226, 8'd228}: color_data = 12'h500;
			{9'd226, 8'd229}: color_data = 12'h500;
			{9'd226, 8'd230}: color_data = 12'h100;
			{9'd226, 8'd231}: color_data = 12'h710;
			{9'd226, 8'd232}: color_data = 12'hc10;
			{9'd226, 8'd233}: color_data = 12'h900;
			{9'd226, 8'd234}: color_data = 12'h500;
			{9'd226, 8'd235}: color_data = 12'h100;
			{9'd226, 8'd236}: color_data = 12'h500;
			{9'd226, 8'd237}: color_data = 12'h600;
			{9'd226, 8'd238}: color_data = 12'h400;
			{9'd226, 8'd239}: color_data = 12'h000;
			{9'd227, 8'd68}: color_data = 12'h057;
			{9'd227, 8'd69}: color_data = 12'h3bd;
			{9'd227, 8'd70}: color_data = 12'h555;
			{9'd227, 8'd71}: color_data = 12'h002;
			{9'd227, 8'd72}: color_data = 12'h005;
			{9'd227, 8'd73}: color_data = 12'h005;
			{9'd227, 8'd74}: color_data = 12'h004;
			{9'd227, 8'd75}: color_data = 12'h025;
			{9'd227, 8'd76}: color_data = 12'h09c;
			{9'd227, 8'd77}: color_data = 12'h034;
			{9'd227, 8'd119}: color_data = 12'h000;
			{9'd227, 8'd120}: color_data = 12'h1ac;
			{9'd227, 8'd121}: color_data = 12'h689;
			{9'd227, 8'd122}: color_data = 12'h212;
			{9'd227, 8'd123}: color_data = 12'h004;
			{9'd227, 8'd124}: color_data = 12'h005;
			{9'd227, 8'd125}: color_data = 12'h005;
			{9'd227, 8'd126}: color_data = 12'h003;
			{9'd227, 8'd127}: color_data = 12'h06a;
			{9'd227, 8'd128}: color_data = 12'h079;
			{9'd227, 8'd129}: color_data = 12'h000;
			{9'd227, 8'd170}: color_data = 12'h000;
			{9'd227, 8'd171}: color_data = 12'h079;
			{9'd227, 8'd172}: color_data = 12'h4bd;
			{9'd227, 8'd173}: color_data = 12'h444;
			{9'd227, 8'd174}: color_data = 12'h002;
			{9'd227, 8'd175}: color_data = 12'h005;
			{9'd227, 8'd176}: color_data = 12'h005;
			{9'd227, 8'd177}: color_data = 12'h004;
			{9'd227, 8'd178}: color_data = 12'h036;
			{9'd227, 8'd179}: color_data = 12'h09c;
			{9'd227, 8'd180}: color_data = 12'h023;
			{9'd227, 8'd222}: color_data = 12'h410;
			{9'd227, 8'd223}: color_data = 12'hd30;
			{9'd227, 8'd224}: color_data = 12'hb00;
			{9'd227, 8'd225}: color_data = 12'h700;
			{9'd227, 8'd226}: color_data = 12'h200;
			{9'd227, 8'd227}: color_data = 12'h700;
			{9'd227, 8'd228}: color_data = 12'hb00;
			{9'd227, 8'd229}: color_data = 12'ha00;
			{9'd227, 8'd230}: color_data = 12'h300;
			{9'd227, 8'd231}: color_data = 12'h820;
			{9'd227, 8'd232}: color_data = 12'hd20;
			{9'd227, 8'd233}: color_data = 12'h900;
			{9'd227, 8'd234}: color_data = 12'h500;
			{9'd227, 8'd235}: color_data = 12'h300;
			{9'd227, 8'd236}: color_data = 12'h900;
			{9'd227, 8'd237}: color_data = 12'hb00;
			{9'd227, 8'd238}: color_data = 12'h800;
			{9'd227, 8'd239}: color_data = 12'h100;
			{9'd228, 8'd68}: color_data = 12'h035;
			{9'd228, 8'd69}: color_data = 12'h047;
			{9'd228, 8'd70}: color_data = 12'h001;
			{9'd228, 8'd71}: color_data = 12'h004;
			{9'd228, 8'd72}: color_data = 12'h004;
			{9'd228, 8'd73}: color_data = 12'h004;
			{9'd228, 8'd74}: color_data = 12'h004;
			{9'd228, 8'd75}: color_data = 12'h015;
			{9'd228, 8'd76}: color_data = 12'h059;
			{9'd228, 8'd77}: color_data = 12'h023;
			{9'd228, 8'd119}: color_data = 12'h000;
			{9'd228, 8'd120}: color_data = 12'h058;
			{9'd228, 8'd121}: color_data = 12'h013;
			{9'd228, 8'd122}: color_data = 12'h002;
			{9'd228, 8'd123}: color_data = 12'h004;
			{9'd228, 8'd124}: color_data = 12'h004;
			{9'd228, 8'd125}: color_data = 12'h004;
			{9'd228, 8'd126}: color_data = 12'h004;
			{9'd228, 8'd127}: color_data = 12'h038;
			{9'd228, 8'd128}: color_data = 12'h046;
			{9'd228, 8'd129}: color_data = 12'h000;
			{9'd228, 8'd170}: color_data = 12'h000;
			{9'd228, 8'd171}: color_data = 12'h047;
			{9'd228, 8'd172}: color_data = 12'h036;
			{9'd228, 8'd173}: color_data = 12'h001;
			{9'd228, 8'd174}: color_data = 12'h004;
			{9'd228, 8'd175}: color_data = 12'h004;
			{9'd228, 8'd176}: color_data = 12'h004;
			{9'd228, 8'd177}: color_data = 12'h004;
			{9'd228, 8'd178}: color_data = 12'h016;
			{9'd228, 8'd179}: color_data = 12'h059;
			{9'd228, 8'd180}: color_data = 12'h012;
			{9'd228, 8'd222}: color_data = 12'h410;
			{9'd228, 8'd223}: color_data = 12'he40;
			{9'd228, 8'd224}: color_data = 12'hd20;
			{9'd228, 8'd225}: color_data = 12'h800;
			{9'd228, 8'd226}: color_data = 12'h200;
			{9'd228, 8'd227}: color_data = 12'h600;
			{9'd228, 8'd228}: color_data = 12'ha00;
			{9'd228, 8'd229}: color_data = 12'h900;
			{9'd228, 8'd230}: color_data = 12'h300;
			{9'd228, 8'd231}: color_data = 12'h820;
			{9'd228, 8'd232}: color_data = 12'hf30;
			{9'd228, 8'd233}: color_data = 12'hc00;
			{9'd228, 8'd234}: color_data = 12'h500;
			{9'd228, 8'd235}: color_data = 12'h200;
			{9'd228, 8'd236}: color_data = 12'h900;
			{9'd228, 8'd237}: color_data = 12'ha00;
			{9'd228, 8'd238}: color_data = 12'h700;
			{9'd228, 8'd239}: color_data = 12'h100;
			{9'd229, 8'd68}: color_data = 12'h013;
			{9'd229, 8'd69}: color_data = 12'h027;
			{9'd229, 8'd70}: color_data = 12'h016;
			{9'd229, 8'd71}: color_data = 12'h027;
			{9'd229, 8'd72}: color_data = 12'h027;
			{9'd229, 8'd73}: color_data = 12'h017;
			{9'd229, 8'd74}: color_data = 12'h027;
			{9'd229, 8'd75}: color_data = 12'h028;
			{9'd229, 8'd76}: color_data = 12'h027;
			{9'd229, 8'd77}: color_data = 12'h001;
			{9'd229, 8'd119}: color_data = 12'h000;
			{9'd229, 8'd120}: color_data = 12'h016;
			{9'd229, 8'd121}: color_data = 12'h017;
			{9'd229, 8'd122}: color_data = 12'h017;
			{9'd229, 8'd123}: color_data = 12'h027;
			{9'd229, 8'd124}: color_data = 12'h027;
			{9'd229, 8'd125}: color_data = 12'h027;
			{9'd229, 8'd126}: color_data = 12'h027;
			{9'd229, 8'd127}: color_data = 12'h028;
			{9'd229, 8'd128}: color_data = 12'h014;
			{9'd229, 8'd129}: color_data = 12'h000;
			{9'd229, 8'd170}: color_data = 12'h000;
			{9'd229, 8'd171}: color_data = 12'h014;
			{9'd229, 8'd172}: color_data = 12'h027;
			{9'd229, 8'd173}: color_data = 12'h016;
			{9'd229, 8'd174}: color_data = 12'h027;
			{9'd229, 8'd175}: color_data = 12'h027;
			{9'd229, 8'd176}: color_data = 12'h027;
			{9'd229, 8'd177}: color_data = 12'h027;
			{9'd229, 8'd178}: color_data = 12'h028;
			{9'd229, 8'd179}: color_data = 12'h026;
			{9'd229, 8'd180}: color_data = 12'h001;
			{9'd229, 8'd222}: color_data = 12'h300;
			{9'd229, 8'd223}: color_data = 12'hc30;
			{9'd229, 8'd224}: color_data = 12'hc30;
			{9'd229, 8'd225}: color_data = 12'h600;
			{9'd229, 8'd226}: color_data = 12'h100;
			{9'd229, 8'd227}: color_data = 12'h600;
			{9'd229, 8'd228}: color_data = 12'ha00;
			{9'd229, 8'd229}: color_data = 12'h900;
			{9'd229, 8'd230}: color_data = 12'h300;
			{9'd229, 8'd231}: color_data = 12'h620;
			{9'd229, 8'd232}: color_data = 12'hd40;
			{9'd229, 8'd233}: color_data = 12'ha20;
			{9'd229, 8'd234}: color_data = 12'h300;
			{9'd229, 8'd235}: color_data = 12'h200;
			{9'd229, 8'd236}: color_data = 12'h900;
			{9'd229, 8'd237}: color_data = 12'ha00;
			{9'd229, 8'd238}: color_data = 12'h700;
			{9'd229, 8'd239}: color_data = 12'h100;
			{9'd230, 8'd68}: color_data = 12'h035;
			{9'd230, 8'd69}: color_data = 12'h09e;
			{9'd230, 8'd70}: color_data = 12'h09e;
			{9'd230, 8'd71}: color_data = 12'h09e;
			{9'd230, 8'd72}: color_data = 12'h09e;
			{9'd230, 8'd73}: color_data = 12'h09e;
			{9'd230, 8'd74}: color_data = 12'h09e;
			{9'd230, 8'd75}: color_data = 12'h09e;
			{9'd230, 8'd76}: color_data = 12'h08c;
			{9'd230, 8'd77}: color_data = 12'h023;
			{9'd230, 8'd119}: color_data = 12'h000;
			{9'd230, 8'd120}: color_data = 12'h07b;
			{9'd230, 8'd121}: color_data = 12'h0ae;
			{9'd230, 8'd122}: color_data = 12'h09e;
			{9'd230, 8'd123}: color_data = 12'h09e;
			{9'd230, 8'd124}: color_data = 12'h09e;
			{9'd230, 8'd125}: color_data = 12'h09e;
			{9'd230, 8'd126}: color_data = 12'h09e;
			{9'd230, 8'd127}: color_data = 12'h09e;
			{9'd230, 8'd128}: color_data = 12'h057;
			{9'd230, 8'd129}: color_data = 12'h000;
			{9'd230, 8'd170}: color_data = 12'h000;
			{9'd230, 8'd171}: color_data = 12'h057;
			{9'd230, 8'd172}: color_data = 12'h0ae;
			{9'd230, 8'd173}: color_data = 12'h09e;
			{9'd230, 8'd174}: color_data = 12'h09e;
			{9'd230, 8'd175}: color_data = 12'h09e;
			{9'd230, 8'd176}: color_data = 12'h09e;
			{9'd230, 8'd177}: color_data = 12'h09e;
			{9'd230, 8'd178}: color_data = 12'h09e;
			{9'd230, 8'd179}: color_data = 12'h07b;
			{9'd230, 8'd180}: color_data = 12'h012;
			{9'd230, 8'd222}: color_data = 12'h000;
			{9'd230, 8'd223}: color_data = 12'h200;
			{9'd230, 8'd224}: color_data = 12'h300;
			{9'd230, 8'd225}: color_data = 12'h100;
			{9'd230, 8'd226}: color_data = 12'h000;
			{9'd230, 8'd227}: color_data = 12'h700;
			{9'd230, 8'd228}: color_data = 12'ha00;
			{9'd230, 8'd229}: color_data = 12'h900;
			{9'd230, 8'd230}: color_data = 12'h300;
			{9'd230, 8'd231}: color_data = 12'h100;
			{9'd230, 8'd232}: color_data = 12'h310;
			{9'd230, 8'd233}: color_data = 12'h200;
			{9'd230, 8'd234}: color_data = 12'h000;
			{9'd230, 8'd235}: color_data = 12'h300;
			{9'd230, 8'd236}: color_data = 12'h900;
			{9'd230, 8'd237}: color_data = 12'ha00;
			{9'd230, 8'd238}: color_data = 12'h700;
			{9'd230, 8'd239}: color_data = 12'h100;
			{9'd231, 8'd68}: color_data = 12'h057;
			{9'd231, 8'd69}: color_data = 12'h4ef;
			{9'd231, 8'd70}: color_data = 12'h7ef;
			{9'd231, 8'd71}: color_data = 12'h0cf;
			{9'd231, 8'd72}: color_data = 12'h0cf;
			{9'd231, 8'd73}: color_data = 12'h0df;
			{9'd231, 8'd74}: color_data = 12'h0bd;
			{9'd231, 8'd75}: color_data = 12'h068;
			{9'd231, 8'd76}: color_data = 12'h09c;
			{9'd231, 8'd77}: color_data = 12'h034;
			{9'd231, 8'd119}: color_data = 12'h000;
			{9'd231, 8'd120}: color_data = 12'h1ad;
			{9'd231, 8'd121}: color_data = 12'h8ff;
			{9'd231, 8'd122}: color_data = 12'h3df;
			{9'd231, 8'd123}: color_data = 12'h0cf;
			{9'd231, 8'd124}: color_data = 12'h0cf;
			{9'd231, 8'd125}: color_data = 12'h0cf;
			{9'd231, 8'd126}: color_data = 12'h07a;
			{9'd231, 8'd127}: color_data = 12'h08b;
			{9'd231, 8'd128}: color_data = 12'h079;
			{9'd231, 8'd129}: color_data = 12'h000;
			{9'd231, 8'd170}: color_data = 12'h000;
			{9'd231, 8'd171}: color_data = 12'h069;
			{9'd231, 8'd172}: color_data = 12'h6ef;
			{9'd231, 8'd173}: color_data = 12'h6ef;
			{9'd231, 8'd174}: color_data = 12'h0cf;
			{9'd231, 8'd175}: color_data = 12'h0cf;
			{9'd231, 8'd176}: color_data = 12'h0df;
			{9'd231, 8'd177}: color_data = 12'h0ac;
			{9'd231, 8'd178}: color_data = 12'h079;
			{9'd231, 8'd179}: color_data = 12'h09c;
			{9'd231, 8'd180}: color_data = 12'h023;
			{9'd231, 8'd222}: color_data = 12'h100;
			{9'd231, 8'd223}: color_data = 12'h400;
			{9'd231, 8'd224}: color_data = 12'h500;
			{9'd231, 8'd225}: color_data = 12'h400;
			{9'd231, 8'd226}: color_data = 12'h200;
			{9'd231, 8'd227}: color_data = 12'ha20;
			{9'd231, 8'd228}: color_data = 12'hb10;
			{9'd231, 8'd229}: color_data = 12'h900;
			{9'd231, 8'd230}: color_data = 12'h300;
			{9'd231, 8'd231}: color_data = 12'h200;
			{9'd231, 8'd232}: color_data = 12'h500;
			{9'd231, 8'd233}: color_data = 12'h500;
			{9'd231, 8'd234}: color_data = 12'h200;
			{9'd231, 8'd235}: color_data = 12'h410;
			{9'd231, 8'd236}: color_data = 12'hc20;
			{9'd231, 8'd237}: color_data = 12'ha00;
			{9'd231, 8'd238}: color_data = 12'h700;
			{9'd231, 8'd239}: color_data = 12'h100;
			{9'd232, 8'd68}: color_data = 12'h047;
			{9'd232, 8'd69}: color_data = 12'h6df;
			{9'd232, 8'd70}: color_data = 12'heff;
			{9'd232, 8'd71}: color_data = 12'h6df;
			{9'd232, 8'd72}: color_data = 12'h0bf;
			{9'd232, 8'd73}: color_data = 12'h0be;
			{9'd232, 8'd74}: color_data = 12'h056;
			{9'd232, 8'd75}: color_data = 12'h012;
			{9'd232, 8'd76}: color_data = 12'h08b;
			{9'd232, 8'd77}: color_data = 12'h034;
			{9'd232, 8'd119}: color_data = 12'h000;
			{9'd232, 8'd120}: color_data = 12'h2ac;
			{9'd232, 8'd121}: color_data = 12'hdff;
			{9'd232, 8'd122}: color_data = 12'haef;
			{9'd232, 8'd123}: color_data = 12'h1bf;
			{9'd232, 8'd124}: color_data = 12'h0cf;
			{9'd232, 8'd125}: color_data = 12'h08b;
			{9'd232, 8'd126}: color_data = 12'h012;
			{9'd232, 8'd127}: color_data = 12'h068;
			{9'd232, 8'd128}: color_data = 12'h079;
			{9'd232, 8'd129}: color_data = 12'h000;
			{9'd232, 8'd170}: color_data = 12'h000;
			{9'd232, 8'd171}: color_data = 12'h068;
			{9'd232, 8'd172}: color_data = 12'h8ef;
			{9'd232, 8'd173}: color_data = 12'hdff;
			{9'd232, 8'd174}: color_data = 12'h4cf;
			{9'd232, 8'd175}: color_data = 12'h0cf;
			{9'd232, 8'd176}: color_data = 12'h0ae;
			{9'd232, 8'd177}: color_data = 12'h035;
			{9'd232, 8'd178}: color_data = 12'h023;
			{9'd232, 8'd179}: color_data = 12'h08c;
			{9'd232, 8'd180}: color_data = 12'h023;
			{9'd232, 8'd222}: color_data = 12'h200;
			{9'd232, 8'd223}: color_data = 12'h900;
			{9'd232, 8'd224}: color_data = 12'hb00;
			{9'd232, 8'd225}: color_data = 12'h800;
			{9'd232, 8'd226}: color_data = 12'h200;
			{9'd232, 8'd227}: color_data = 12'hb30;
			{9'd232, 8'd228}: color_data = 12'hc10;
			{9'd232, 8'd229}: color_data = 12'h800;
			{9'd232, 8'd230}: color_data = 12'h300;
			{9'd232, 8'd231}: color_data = 12'h400;
			{9'd232, 8'd232}: color_data = 12'ha00;
			{9'd232, 8'd233}: color_data = 12'ha00;
			{9'd232, 8'd234}: color_data = 12'h500;
			{9'd232, 8'd235}: color_data = 12'h510;
			{9'd232, 8'd236}: color_data = 12'hd30;
			{9'd232, 8'd237}: color_data = 12'ha00;
			{9'd232, 8'd238}: color_data = 12'h700;
			{9'd232, 8'd239}: color_data = 12'h100;
			{9'd233, 8'd68}: color_data = 12'h047;
			{9'd233, 8'd69}: color_data = 12'h6df;
			{9'd233, 8'd70}: color_data = 12'hfff;
			{9'd233, 8'd71}: color_data = 12'hdff;
			{9'd233, 8'd72}: color_data = 12'h5df;
			{9'd233, 8'd73}: color_data = 12'h068;
			{9'd233, 8'd74}: color_data = 12'h000;
			{9'd233, 8'd75}: color_data = 12'h012;
			{9'd233, 8'd76}: color_data = 12'h08c;
			{9'd233, 8'd77}: color_data = 12'h034;
			{9'd233, 8'd119}: color_data = 12'h000;
			{9'd233, 8'd120}: color_data = 12'h1ac;
			{9'd233, 8'd121}: color_data = 12'hdff;
			{9'd233, 8'd122}: color_data = 12'hfff;
			{9'd233, 8'd123}: color_data = 12'h8ef;
			{9'd233, 8'd124}: color_data = 12'h19c;
			{9'd233, 8'd125}: color_data = 12'h023;
			{9'd233, 8'd127}: color_data = 12'h068;
			{9'd233, 8'd128}: color_data = 12'h079;
			{9'd233, 8'd129}: color_data = 12'h000;
			{9'd233, 8'd170}: color_data = 12'h000;
			{9'd233, 8'd171}: color_data = 12'h068;
			{9'd233, 8'd172}: color_data = 12'h8ef;
			{9'd233, 8'd173}: color_data = 12'hfff;
			{9'd233, 8'd174}: color_data = 12'hcff;
			{9'd233, 8'd175}: color_data = 12'h4ce;
			{9'd233, 8'd176}: color_data = 12'h057;
			{9'd233, 8'd177}: color_data = 12'h000;
			{9'd233, 8'd178}: color_data = 12'h023;
			{9'd233, 8'd179}: color_data = 12'h08c;
			{9'd233, 8'd180}: color_data = 12'h023;
			{9'd233, 8'd222}: color_data = 12'h200;
			{9'd233, 8'd223}: color_data = 12'h900;
			{9'd233, 8'd224}: color_data = 12'ha00;
			{9'd233, 8'd225}: color_data = 12'h700;
			{9'd233, 8'd226}: color_data = 12'h200;
			{9'd233, 8'd227}: color_data = 12'hb30;
			{9'd233, 8'd228}: color_data = 12'he20;
			{9'd233, 8'd229}: color_data = 12'ha00;
			{9'd233, 8'd230}: color_data = 12'h300;
			{9'd233, 8'd231}: color_data = 12'h400;
			{9'd233, 8'd232}: color_data = 12'ha00;
			{9'd233, 8'd233}: color_data = 12'ha00;
			{9'd233, 8'd234}: color_data = 12'h400;
			{9'd233, 8'd235}: color_data = 12'h510;
			{9'd233, 8'd236}: color_data = 12'hf40;
			{9'd233, 8'd237}: color_data = 12'hd10;
			{9'd233, 8'd238}: color_data = 12'h800;
			{9'd233, 8'd239}: color_data = 12'h100;
			{9'd234, 8'd68}: color_data = 12'h047;
			{9'd234, 8'd69}: color_data = 12'h6df;
			{9'd234, 8'd70}: color_data = 12'hfff;
			{9'd234, 8'd71}: color_data = 12'hfff;
			{9'd234, 8'd72}: color_data = 12'h9aa;
			{9'd234, 8'd73}: color_data = 12'h011;
			{9'd234, 8'd75}: color_data = 12'h012;
			{9'd234, 8'd76}: color_data = 12'h08c;
			{9'd234, 8'd77}: color_data = 12'h034;
			{9'd234, 8'd119}: color_data = 12'h000;
			{9'd234, 8'd120}: color_data = 12'h1ac;
			{9'd234, 8'd121}: color_data = 12'hcff;
			{9'd234, 8'd122}: color_data = 12'hfff;
			{9'd234, 8'd123}: color_data = 12'hddd;
			{9'd234, 8'd124}: color_data = 12'h345;
			{9'd234, 8'd126}: color_data = 12'h000;
			{9'd234, 8'd127}: color_data = 12'h068;
			{9'd234, 8'd128}: color_data = 12'h079;
			{9'd234, 8'd129}: color_data = 12'h000;
			{9'd234, 8'd170}: color_data = 12'h000;
			{9'd234, 8'd171}: color_data = 12'h068;
			{9'd234, 8'd172}: color_data = 12'h7ef;
			{9'd234, 8'd173}: color_data = 12'hfff;
			{9'd234, 8'd174}: color_data = 12'hfff;
			{9'd234, 8'd175}: color_data = 12'h899;
			{9'd234, 8'd176}: color_data = 12'h001;
			{9'd234, 8'd178}: color_data = 12'h024;
			{9'd234, 8'd179}: color_data = 12'h08c;
			{9'd234, 8'd180}: color_data = 12'h023;
			{9'd234, 8'd222}: color_data = 12'h200;
			{9'd234, 8'd223}: color_data = 12'h800;
			{9'd234, 8'd224}: color_data = 12'ha00;
			{9'd234, 8'd225}: color_data = 12'h700;
			{9'd234, 8'd226}: color_data = 12'h200;
			{9'd234, 8'd227}: color_data = 12'h920;
			{9'd234, 8'd228}: color_data = 12'hd30;
			{9'd234, 8'd229}: color_data = 12'h910;
			{9'd234, 8'd230}: color_data = 12'h200;
			{9'd234, 8'd231}: color_data = 12'h400;
			{9'd234, 8'd232}: color_data = 12'h900;
			{9'd234, 8'd233}: color_data = 12'ha00;
			{9'd234, 8'd234}: color_data = 12'h400;
			{9'd234, 8'd235}: color_data = 12'h310;
			{9'd234, 8'd236}: color_data = 12'hc30;
			{9'd234, 8'd237}: color_data = 12'hc20;
			{9'd234, 8'd238}: color_data = 12'h600;
			{9'd234, 8'd239}: color_data = 12'h000;
			{9'd235, 8'd68}: color_data = 12'h047;
			{9'd235, 8'd69}: color_data = 12'h6df;
			{9'd235, 8'd70}: color_data = 12'hfff;
			{9'd235, 8'd71}: color_data = 12'hcbb;
			{9'd235, 8'd72}: color_data = 12'h323;
			{9'd235, 8'd73}: color_data = 12'h002;
			{9'd235, 8'd74}: color_data = 12'h000;
			{9'd235, 8'd75}: color_data = 12'h012;
			{9'd235, 8'd76}: color_data = 12'h08c;
			{9'd235, 8'd77}: color_data = 12'h034;
			{9'd235, 8'd119}: color_data = 12'h000;
			{9'd235, 8'd120}: color_data = 12'h1ac;
			{9'd235, 8'd121}: color_data = 12'hdff;
			{9'd235, 8'd122}: color_data = 12'hfee;
			{9'd235, 8'd123}: color_data = 12'h666;
			{9'd235, 8'd124}: color_data = 12'h002;
			{9'd235, 8'd125}: color_data = 12'h001;
			{9'd235, 8'd126}: color_data = 12'h000;
			{9'd235, 8'd127}: color_data = 12'h068;
			{9'd235, 8'd128}: color_data = 12'h079;
			{9'd235, 8'd129}: color_data = 12'h000;
			{9'd235, 8'd170}: color_data = 12'h000;
			{9'd235, 8'd171}: color_data = 12'h068;
			{9'd235, 8'd172}: color_data = 12'h8ef;
			{9'd235, 8'd173}: color_data = 12'hfff;
			{9'd235, 8'd174}: color_data = 12'haa9;
			{9'd235, 8'd175}: color_data = 12'h212;
			{9'd235, 8'd176}: color_data = 12'h002;
			{9'd235, 8'd178}: color_data = 12'h023;
			{9'd235, 8'd179}: color_data = 12'h08c;
			{9'd235, 8'd180}: color_data = 12'h023;
			{9'd235, 8'd222}: color_data = 12'h200;
			{9'd235, 8'd223}: color_data = 12'h900;
			{9'd235, 8'd224}: color_data = 12'ha00;
			{9'd235, 8'd225}: color_data = 12'h800;
			{9'd235, 8'd226}: color_data = 12'h100;
			{9'd235, 8'd227}: color_data = 12'h100;
			{9'd235, 8'd228}: color_data = 12'h310;
			{9'd235, 8'd229}: color_data = 12'h200;
			{9'd235, 8'd230}: color_data = 12'h000;
			{9'd235, 8'd231}: color_data = 12'h500;
			{9'd235, 8'd232}: color_data = 12'ha00;
			{9'd235, 8'd233}: color_data = 12'ha00;
			{9'd235, 8'd234}: color_data = 12'h500;
			{9'd235, 8'd235}: color_data = 12'h000;
			{9'd235, 8'd236}: color_data = 12'h200;
			{9'd235, 8'd237}: color_data = 12'h300;
			{9'd235, 8'd238}: color_data = 12'h100;
			{9'd235, 8'd239}: color_data = 12'h000;
			{9'd236, 8'd68}: color_data = 12'h047;
			{9'd236, 8'd69}: color_data = 12'h6ef;
			{9'd236, 8'd70}: color_data = 12'hdcc;
			{9'd236, 8'd71}: color_data = 12'h434;
			{9'd236, 8'd72}: color_data = 12'h003;
			{9'd236, 8'd73}: color_data = 12'h005;
			{9'd236, 8'd74}: color_data = 12'h002;
			{9'd236, 8'd75}: color_data = 12'h012;
			{9'd236, 8'd76}: color_data = 12'h08c;
			{9'd236, 8'd77}: color_data = 12'h034;
			{9'd236, 8'd119}: color_data = 12'h000;
			{9'd236, 8'd120}: color_data = 12'h2ad;
			{9'd236, 8'd121}: color_data = 12'hcff;
			{9'd236, 8'd122}: color_data = 12'h877;
			{9'd236, 8'd123}: color_data = 12'h002;
			{9'd236, 8'd124}: color_data = 12'h004;
			{9'd236, 8'd125}: color_data = 12'h004;
			{9'd236, 8'd126}: color_data = 12'h000;
			{9'd236, 8'd127}: color_data = 12'h068;
			{9'd236, 8'd128}: color_data = 12'h079;
			{9'd236, 8'd129}: color_data = 12'h000;
			{9'd236, 8'd170}: color_data = 12'h000;
			{9'd236, 8'd171}: color_data = 12'h068;
			{9'd236, 8'd172}: color_data = 12'h8ff;
			{9'd236, 8'd173}: color_data = 12'hcbb;
			{9'd236, 8'd174}: color_data = 12'h223;
			{9'd236, 8'd175}: color_data = 12'h003;
			{9'd236, 8'd176}: color_data = 12'h005;
			{9'd236, 8'd177}: color_data = 12'h002;
			{9'd236, 8'd178}: color_data = 12'h023;
			{9'd236, 8'd179}: color_data = 12'h09c;
			{9'd236, 8'd180}: color_data = 12'h023;
			{9'd236, 8'd222}: color_data = 12'h300;
			{9'd236, 8'd223}: color_data = 12'hc20;
			{9'd236, 8'd224}: color_data = 12'ha00;
			{9'd236, 8'd225}: color_data = 12'h800;
			{9'd236, 8'd226}: color_data = 12'h100;
			{9'd236, 8'd227}: color_data = 12'h300;
			{9'd236, 8'd228}: color_data = 12'h500;
			{9'd236, 8'd229}: color_data = 12'h500;
			{9'd236, 8'd230}: color_data = 12'h100;
			{9'd236, 8'd231}: color_data = 12'h710;
			{9'd236, 8'd232}: color_data = 12'hc10;
			{9'd236, 8'd233}: color_data = 12'h900;
			{9'd236, 8'd234}: color_data = 12'h500;
			{9'd236, 8'd235}: color_data = 12'h100;
			{9'd236, 8'd236}: color_data = 12'h500;
			{9'd236, 8'd237}: color_data = 12'h600;
			{9'd236, 8'd238}: color_data = 12'h400;
			{9'd236, 8'd239}: color_data = 12'h000;
			{9'd237, 8'd68}: color_data = 12'h057;
			{9'd237, 8'd69}: color_data = 12'h3bd;
			{9'd237, 8'd70}: color_data = 12'h555;
			{9'd237, 8'd71}: color_data = 12'h002;
			{9'd237, 8'd72}: color_data = 12'h005;
			{9'd237, 8'd73}: color_data = 12'h005;
			{9'd237, 8'd74}: color_data = 12'h004;
			{9'd237, 8'd75}: color_data = 12'h025;
			{9'd237, 8'd76}: color_data = 12'h09c;
			{9'd237, 8'd77}: color_data = 12'h034;
			{9'd237, 8'd119}: color_data = 12'h000;
			{9'd237, 8'd120}: color_data = 12'h1ac;
			{9'd237, 8'd121}: color_data = 12'h689;
			{9'd237, 8'd122}: color_data = 12'h212;
			{9'd237, 8'd123}: color_data = 12'h004;
			{9'd237, 8'd124}: color_data = 12'h005;
			{9'd237, 8'd125}: color_data = 12'h005;
			{9'd237, 8'd126}: color_data = 12'h003;
			{9'd237, 8'd127}: color_data = 12'h06a;
			{9'd237, 8'd128}: color_data = 12'h079;
			{9'd237, 8'd129}: color_data = 12'h000;
			{9'd237, 8'd170}: color_data = 12'h000;
			{9'd237, 8'd171}: color_data = 12'h079;
			{9'd237, 8'd172}: color_data = 12'h4bd;
			{9'd237, 8'd173}: color_data = 12'h444;
			{9'd237, 8'd174}: color_data = 12'h002;
			{9'd237, 8'd175}: color_data = 12'h005;
			{9'd237, 8'd176}: color_data = 12'h005;
			{9'd237, 8'd177}: color_data = 12'h004;
			{9'd237, 8'd178}: color_data = 12'h036;
			{9'd237, 8'd179}: color_data = 12'h09c;
			{9'd237, 8'd180}: color_data = 12'h023;
			{9'd237, 8'd222}: color_data = 12'h410;
			{9'd237, 8'd223}: color_data = 12'hd30;
			{9'd237, 8'd224}: color_data = 12'hb00;
			{9'd237, 8'd225}: color_data = 12'h700;
			{9'd237, 8'd226}: color_data = 12'h200;
			{9'd237, 8'd227}: color_data = 12'h700;
			{9'd237, 8'd228}: color_data = 12'hb00;
			{9'd237, 8'd229}: color_data = 12'ha00;
			{9'd237, 8'd230}: color_data = 12'h300;
			{9'd237, 8'd231}: color_data = 12'h820;
			{9'd237, 8'd232}: color_data = 12'hd20;
			{9'd237, 8'd233}: color_data = 12'h900;
			{9'd237, 8'd234}: color_data = 12'h500;
			{9'd237, 8'd235}: color_data = 12'h300;
			{9'd237, 8'd236}: color_data = 12'h900;
			{9'd237, 8'd237}: color_data = 12'hb00;
			{9'd237, 8'd238}: color_data = 12'h800;
			{9'd237, 8'd239}: color_data = 12'h100;
			{9'd238, 8'd68}: color_data = 12'h035;
			{9'd238, 8'd69}: color_data = 12'h047;
			{9'd238, 8'd70}: color_data = 12'h001;
			{9'd238, 8'd71}: color_data = 12'h004;
			{9'd238, 8'd72}: color_data = 12'h004;
			{9'd238, 8'd73}: color_data = 12'h004;
			{9'd238, 8'd74}: color_data = 12'h004;
			{9'd238, 8'd75}: color_data = 12'h015;
			{9'd238, 8'd76}: color_data = 12'h059;
			{9'd238, 8'd77}: color_data = 12'h023;
			{9'd238, 8'd119}: color_data = 12'h000;
			{9'd238, 8'd120}: color_data = 12'h058;
			{9'd238, 8'd121}: color_data = 12'h013;
			{9'd238, 8'd122}: color_data = 12'h002;
			{9'd238, 8'd123}: color_data = 12'h004;
			{9'd238, 8'd124}: color_data = 12'h004;
			{9'd238, 8'd125}: color_data = 12'h004;
			{9'd238, 8'd126}: color_data = 12'h004;
			{9'd238, 8'd127}: color_data = 12'h038;
			{9'd238, 8'd128}: color_data = 12'h046;
			{9'd238, 8'd129}: color_data = 12'h000;
			{9'd238, 8'd170}: color_data = 12'h000;
			{9'd238, 8'd171}: color_data = 12'h047;
			{9'd238, 8'd172}: color_data = 12'h036;
			{9'd238, 8'd173}: color_data = 12'h001;
			{9'd238, 8'd174}: color_data = 12'h004;
			{9'd238, 8'd175}: color_data = 12'h004;
			{9'd238, 8'd176}: color_data = 12'h004;
			{9'd238, 8'd177}: color_data = 12'h004;
			{9'd238, 8'd178}: color_data = 12'h016;
			{9'd238, 8'd179}: color_data = 12'h059;
			{9'd238, 8'd180}: color_data = 12'h012;
			{9'd238, 8'd222}: color_data = 12'h410;
			{9'd238, 8'd223}: color_data = 12'he40;
			{9'd238, 8'd224}: color_data = 12'hd20;
			{9'd238, 8'd225}: color_data = 12'h800;
			{9'd238, 8'd226}: color_data = 12'h200;
			{9'd238, 8'd227}: color_data = 12'h600;
			{9'd238, 8'd228}: color_data = 12'ha00;
			{9'd238, 8'd229}: color_data = 12'h900;
			{9'd238, 8'd230}: color_data = 12'h300;
			{9'd238, 8'd231}: color_data = 12'h820;
			{9'd238, 8'd232}: color_data = 12'hf30;
			{9'd238, 8'd233}: color_data = 12'hc00;
			{9'd238, 8'd234}: color_data = 12'h500;
			{9'd238, 8'd235}: color_data = 12'h200;
			{9'd238, 8'd236}: color_data = 12'h900;
			{9'd238, 8'd237}: color_data = 12'ha00;
			{9'd238, 8'd238}: color_data = 12'h700;
			{9'd238, 8'd239}: color_data = 12'h100;
			{9'd239, 8'd68}: color_data = 12'h013;
			{9'd239, 8'd69}: color_data = 12'h027;
			{9'd239, 8'd70}: color_data = 12'h016;
			{9'd239, 8'd71}: color_data = 12'h027;
			{9'd239, 8'd72}: color_data = 12'h027;
			{9'd239, 8'd73}: color_data = 12'h027;
			{9'd239, 8'd74}: color_data = 12'h027;
			{9'd239, 8'd75}: color_data = 12'h028;
			{9'd239, 8'd76}: color_data = 12'h027;
			{9'd239, 8'd77}: color_data = 12'h001;
			{9'd239, 8'd119}: color_data = 12'h000;
			{9'd239, 8'd120}: color_data = 12'h016;
			{9'd239, 8'd121}: color_data = 12'h017;
			{9'd239, 8'd122}: color_data = 12'h027;
			{9'd239, 8'd123}: color_data = 12'h027;
			{9'd239, 8'd124}: color_data = 12'h027;
			{9'd239, 8'd125}: color_data = 12'h027;
			{9'd239, 8'd126}: color_data = 12'h027;
			{9'd239, 8'd127}: color_data = 12'h028;
			{9'd239, 8'd128}: color_data = 12'h014;
			{9'd239, 8'd129}: color_data = 12'h000;
			{9'd239, 8'd170}: color_data = 12'h000;
			{9'd239, 8'd171}: color_data = 12'h014;
			{9'd239, 8'd172}: color_data = 12'h027;
			{9'd239, 8'd173}: color_data = 12'h016;
			{9'd239, 8'd174}: color_data = 12'h027;
			{9'd239, 8'd175}: color_data = 12'h027;
			{9'd239, 8'd176}: color_data = 12'h027;
			{9'd239, 8'd177}: color_data = 12'h027;
			{9'd239, 8'd178}: color_data = 12'h028;
			{9'd239, 8'd179}: color_data = 12'h026;
			{9'd239, 8'd180}: color_data = 12'h001;
			{9'd239, 8'd222}: color_data = 12'h300;
			{9'd239, 8'd223}: color_data = 12'hc30;
			{9'd239, 8'd224}: color_data = 12'hc30;
			{9'd239, 8'd225}: color_data = 12'h600;
			{9'd239, 8'd226}: color_data = 12'h100;
			{9'd239, 8'd227}: color_data = 12'h600;
			{9'd239, 8'd228}: color_data = 12'ha00;
			{9'd239, 8'd229}: color_data = 12'h900;
			{9'd239, 8'd230}: color_data = 12'h300;
			{9'd239, 8'd231}: color_data = 12'h620;
			{9'd239, 8'd232}: color_data = 12'hd40;
			{9'd239, 8'd233}: color_data = 12'ha20;
			{9'd239, 8'd234}: color_data = 12'h300;
			{9'd239, 8'd235}: color_data = 12'h200;
			{9'd239, 8'd236}: color_data = 12'h900;
			{9'd239, 8'd237}: color_data = 12'ha00;
			{9'd239, 8'd238}: color_data = 12'h700;
			{9'd239, 8'd239}: color_data = 12'h100;
			{9'd240, 8'd68}: color_data = 12'h035;
			{9'd240, 8'd69}: color_data = 12'h09e;
			{9'd240, 8'd70}: color_data = 12'h09e;
			{9'd240, 8'd71}: color_data = 12'h09e;
			{9'd240, 8'd72}: color_data = 12'h09e;
			{9'd240, 8'd73}: color_data = 12'h09e;
			{9'd240, 8'd74}: color_data = 12'h09e;
			{9'd240, 8'd75}: color_data = 12'h09e;
			{9'd240, 8'd76}: color_data = 12'h08c;
			{9'd240, 8'd77}: color_data = 12'h023;
			{9'd240, 8'd119}: color_data = 12'h000;
			{9'd240, 8'd120}: color_data = 12'h07b;
			{9'd240, 8'd121}: color_data = 12'h0ae;
			{9'd240, 8'd122}: color_data = 12'h09e;
			{9'd240, 8'd123}: color_data = 12'h09e;
			{9'd240, 8'd124}: color_data = 12'h09e;
			{9'd240, 8'd125}: color_data = 12'h09e;
			{9'd240, 8'd126}: color_data = 12'h09e;
			{9'd240, 8'd127}: color_data = 12'h09e;
			{9'd240, 8'd128}: color_data = 12'h057;
			{9'd240, 8'd129}: color_data = 12'h000;
			{9'd240, 8'd170}: color_data = 12'h000;
			{9'd240, 8'd171}: color_data = 12'h057;
			{9'd240, 8'd172}: color_data = 12'h0ae;
			{9'd240, 8'd173}: color_data = 12'h09e;
			{9'd240, 8'd174}: color_data = 12'h09e;
			{9'd240, 8'd175}: color_data = 12'h09e;
			{9'd240, 8'd176}: color_data = 12'h09e;
			{9'd240, 8'd177}: color_data = 12'h09e;
			{9'd240, 8'd178}: color_data = 12'h09e;
			{9'd240, 8'd179}: color_data = 12'h07b;
			{9'd240, 8'd180}: color_data = 12'h012;
			{9'd240, 8'd222}: color_data = 12'h000;
			{9'd240, 8'd223}: color_data = 12'h200;
			{9'd240, 8'd224}: color_data = 12'h300;
			{9'd240, 8'd225}: color_data = 12'h100;
			{9'd240, 8'd226}: color_data = 12'h000;
			{9'd240, 8'd227}: color_data = 12'h700;
			{9'd240, 8'd228}: color_data = 12'ha00;
			{9'd240, 8'd229}: color_data = 12'h900;
			{9'd240, 8'd230}: color_data = 12'h300;
			{9'd240, 8'd231}: color_data = 12'h100;
			{9'd240, 8'd232}: color_data = 12'h300;
			{9'd240, 8'd233}: color_data = 12'h200;
			{9'd240, 8'd234}: color_data = 12'h000;
			{9'd240, 8'd235}: color_data = 12'h300;
			{9'd240, 8'd236}: color_data = 12'h900;
			{9'd240, 8'd237}: color_data = 12'ha00;
			{9'd240, 8'd238}: color_data = 12'h700;
			{9'd240, 8'd239}: color_data = 12'h100;
			{9'd241, 8'd68}: color_data = 12'h057;
			{9'd241, 8'd69}: color_data = 12'h4ef;
			{9'd241, 8'd70}: color_data = 12'h7ef;
			{9'd241, 8'd71}: color_data = 12'h0cf;
			{9'd241, 8'd72}: color_data = 12'h0cf;
			{9'd241, 8'd73}: color_data = 12'h0df;
			{9'd241, 8'd74}: color_data = 12'h0bd;
			{9'd241, 8'd75}: color_data = 12'h068;
			{9'd241, 8'd76}: color_data = 12'h09c;
			{9'd241, 8'd77}: color_data = 12'h034;
			{9'd241, 8'd119}: color_data = 12'h000;
			{9'd241, 8'd120}: color_data = 12'h1ad;
			{9'd241, 8'd121}: color_data = 12'h8ff;
			{9'd241, 8'd122}: color_data = 12'h3df;
			{9'd241, 8'd123}: color_data = 12'h0cf;
			{9'd241, 8'd124}: color_data = 12'h0cf;
			{9'd241, 8'd125}: color_data = 12'h0cf;
			{9'd241, 8'd126}: color_data = 12'h079;
			{9'd241, 8'd127}: color_data = 12'h08b;
			{9'd241, 8'd128}: color_data = 12'h079;
			{9'd241, 8'd129}: color_data = 12'h000;
			{9'd241, 8'd170}: color_data = 12'h000;
			{9'd241, 8'd171}: color_data = 12'h069;
			{9'd241, 8'd172}: color_data = 12'h6ef;
			{9'd241, 8'd173}: color_data = 12'h6ef;
			{9'd241, 8'd174}: color_data = 12'h0cf;
			{9'd241, 8'd175}: color_data = 12'h0cf;
			{9'd241, 8'd176}: color_data = 12'h0df;
			{9'd241, 8'd177}: color_data = 12'h0ac;
			{9'd241, 8'd178}: color_data = 12'h079;
			{9'd241, 8'd179}: color_data = 12'h09c;
			{9'd241, 8'd180}: color_data = 12'h023;
			{9'd241, 8'd222}: color_data = 12'h100;
			{9'd241, 8'd223}: color_data = 12'h500;
			{9'd241, 8'd224}: color_data = 12'h500;
			{9'd241, 8'd225}: color_data = 12'h400;
			{9'd241, 8'd226}: color_data = 12'h200;
			{9'd241, 8'd227}: color_data = 12'ha20;
			{9'd241, 8'd228}: color_data = 12'hb10;
			{9'd241, 8'd229}: color_data = 12'h900;
			{9'd241, 8'd230}: color_data = 12'h300;
			{9'd241, 8'd231}: color_data = 12'h200;
			{9'd241, 8'd232}: color_data = 12'h500;
			{9'd241, 8'd233}: color_data = 12'h500;
			{9'd241, 8'd234}: color_data = 12'h200;
			{9'd241, 8'd235}: color_data = 12'h410;
			{9'd241, 8'd236}: color_data = 12'hc20;
			{9'd241, 8'd237}: color_data = 12'ha00;
			{9'd241, 8'd238}: color_data = 12'h700;
			{9'd241, 8'd239}: color_data = 12'h100;
			{9'd242, 8'd68}: color_data = 12'h047;
			{9'd242, 8'd69}: color_data = 12'h6df;
			{9'd242, 8'd70}: color_data = 12'heff;
			{9'd242, 8'd71}: color_data = 12'h6df;
			{9'd242, 8'd72}: color_data = 12'h0bf;
			{9'd242, 8'd73}: color_data = 12'h0bf;
			{9'd242, 8'd74}: color_data = 12'h056;
			{9'd242, 8'd75}: color_data = 12'h012;
			{9'd242, 8'd76}: color_data = 12'h08b;
			{9'd242, 8'd77}: color_data = 12'h034;
			{9'd242, 8'd119}: color_data = 12'h000;
			{9'd242, 8'd120}: color_data = 12'h2ac;
			{9'd242, 8'd121}: color_data = 12'hdff;
			{9'd242, 8'd122}: color_data = 12'haef;
			{9'd242, 8'd123}: color_data = 12'h1bf;
			{9'd242, 8'd124}: color_data = 12'h0cf;
			{9'd242, 8'd125}: color_data = 12'h08b;
			{9'd242, 8'd126}: color_data = 12'h012;
			{9'd242, 8'd127}: color_data = 12'h068;
			{9'd242, 8'd128}: color_data = 12'h079;
			{9'd242, 8'd129}: color_data = 12'h000;
			{9'd242, 8'd170}: color_data = 12'h000;
			{9'd242, 8'd171}: color_data = 12'h068;
			{9'd242, 8'd172}: color_data = 12'h8ef;
			{9'd242, 8'd173}: color_data = 12'hdff;
			{9'd242, 8'd174}: color_data = 12'h4cf;
			{9'd242, 8'd175}: color_data = 12'h0bf;
			{9'd242, 8'd176}: color_data = 12'h0ae;
			{9'd242, 8'd177}: color_data = 12'h035;
			{9'd242, 8'd178}: color_data = 12'h023;
			{9'd242, 8'd179}: color_data = 12'h08c;
			{9'd242, 8'd180}: color_data = 12'h023;
			{9'd242, 8'd222}: color_data = 12'h200;
			{9'd242, 8'd223}: color_data = 12'h900;
			{9'd242, 8'd224}: color_data = 12'hb00;
			{9'd242, 8'd225}: color_data = 12'h800;
			{9'd242, 8'd226}: color_data = 12'h200;
			{9'd242, 8'd227}: color_data = 12'hb30;
			{9'd242, 8'd228}: color_data = 12'hc10;
			{9'd242, 8'd229}: color_data = 12'h800;
			{9'd242, 8'd230}: color_data = 12'h300;
			{9'd242, 8'd231}: color_data = 12'h400;
			{9'd242, 8'd232}: color_data = 12'ha00;
			{9'd242, 8'd233}: color_data = 12'ha00;
			{9'd242, 8'd234}: color_data = 12'h500;
			{9'd242, 8'd235}: color_data = 12'h510;
			{9'd242, 8'd236}: color_data = 12'hd30;
			{9'd242, 8'd237}: color_data = 12'ha00;
			{9'd242, 8'd238}: color_data = 12'h700;
			{9'd242, 8'd239}: color_data = 12'h100;
			{9'd243, 8'd68}: color_data = 12'h047;
			{9'd243, 8'd69}: color_data = 12'h6df;
			{9'd243, 8'd70}: color_data = 12'hfff;
			{9'd243, 8'd71}: color_data = 12'hdff;
			{9'd243, 8'd72}: color_data = 12'h5df;
			{9'd243, 8'd73}: color_data = 12'h068;
			{9'd243, 8'd74}: color_data = 12'h000;
			{9'd243, 8'd75}: color_data = 12'h012;
			{9'd243, 8'd76}: color_data = 12'h08c;
			{9'd243, 8'd77}: color_data = 12'h034;
			{9'd243, 8'd119}: color_data = 12'h000;
			{9'd243, 8'd120}: color_data = 12'h1ac;
			{9'd243, 8'd121}: color_data = 12'hdff;
			{9'd243, 8'd122}: color_data = 12'hfff;
			{9'd243, 8'd123}: color_data = 12'h9ef;
			{9'd243, 8'd124}: color_data = 12'h19c;
			{9'd243, 8'd125}: color_data = 12'h023;
			{9'd243, 8'd127}: color_data = 12'h068;
			{9'd243, 8'd128}: color_data = 12'h079;
			{9'd243, 8'd129}: color_data = 12'h000;
			{9'd243, 8'd170}: color_data = 12'h000;
			{9'd243, 8'd171}: color_data = 12'h068;
			{9'd243, 8'd172}: color_data = 12'h8ef;
			{9'd243, 8'd173}: color_data = 12'hfff;
			{9'd243, 8'd174}: color_data = 12'hcff;
			{9'd243, 8'd175}: color_data = 12'h4ce;
			{9'd243, 8'd176}: color_data = 12'h057;
			{9'd243, 8'd177}: color_data = 12'h000;
			{9'd243, 8'd178}: color_data = 12'h023;
			{9'd243, 8'd179}: color_data = 12'h08c;
			{9'd243, 8'd180}: color_data = 12'h023;
			{9'd243, 8'd222}: color_data = 12'h200;
			{9'd243, 8'd223}: color_data = 12'h900;
			{9'd243, 8'd224}: color_data = 12'ha00;
			{9'd243, 8'd225}: color_data = 12'h700;
			{9'd243, 8'd226}: color_data = 12'h200;
			{9'd243, 8'd227}: color_data = 12'hb30;
			{9'd243, 8'd228}: color_data = 12'he20;
			{9'd243, 8'd229}: color_data = 12'ha00;
			{9'd243, 8'd230}: color_data = 12'h300;
			{9'd243, 8'd231}: color_data = 12'h400;
			{9'd243, 8'd232}: color_data = 12'ha00;
			{9'd243, 8'd233}: color_data = 12'ha00;
			{9'd243, 8'd234}: color_data = 12'h400;
			{9'd243, 8'd235}: color_data = 12'h510;
			{9'd243, 8'd236}: color_data = 12'hf40;
			{9'd243, 8'd237}: color_data = 12'hd10;
			{9'd243, 8'd238}: color_data = 12'h800;
			{9'd243, 8'd239}: color_data = 12'h100;
			{9'd244, 8'd68}: color_data = 12'h047;
			{9'd244, 8'd69}: color_data = 12'h6df;
			{9'd244, 8'd70}: color_data = 12'hfff;
			{9'd244, 8'd71}: color_data = 12'hfff;
			{9'd244, 8'd72}: color_data = 12'h9aa;
			{9'd244, 8'd73}: color_data = 12'h011;
			{9'd244, 8'd75}: color_data = 12'h012;
			{9'd244, 8'd76}: color_data = 12'h08c;
			{9'd244, 8'd77}: color_data = 12'h034;
			{9'd244, 8'd119}: color_data = 12'h000;
			{9'd244, 8'd120}: color_data = 12'h1ac;
			{9'd244, 8'd121}: color_data = 12'hcff;
			{9'd244, 8'd122}: color_data = 12'hfff;
			{9'd244, 8'd123}: color_data = 12'hddd;
			{9'd244, 8'd124}: color_data = 12'h345;
			{9'd244, 8'd126}: color_data = 12'h000;
			{9'd244, 8'd127}: color_data = 12'h068;
			{9'd244, 8'd128}: color_data = 12'h079;
			{9'd244, 8'd129}: color_data = 12'h000;
			{9'd244, 8'd170}: color_data = 12'h000;
			{9'd244, 8'd171}: color_data = 12'h068;
			{9'd244, 8'd172}: color_data = 12'h7ef;
			{9'd244, 8'd173}: color_data = 12'hfff;
			{9'd244, 8'd174}: color_data = 12'hfff;
			{9'd244, 8'd175}: color_data = 12'h899;
			{9'd244, 8'd176}: color_data = 12'h001;
			{9'd244, 8'd178}: color_data = 12'h024;
			{9'd244, 8'd179}: color_data = 12'h08c;
			{9'd244, 8'd180}: color_data = 12'h023;
			{9'd244, 8'd222}: color_data = 12'h200;
			{9'd244, 8'd223}: color_data = 12'h800;
			{9'd244, 8'd224}: color_data = 12'ha00;
			{9'd244, 8'd225}: color_data = 12'h800;
			{9'd244, 8'd226}: color_data = 12'h200;
			{9'd244, 8'd227}: color_data = 12'h930;
			{9'd244, 8'd228}: color_data = 12'hd30;
			{9'd244, 8'd229}: color_data = 12'h910;
			{9'd244, 8'd230}: color_data = 12'h200;
			{9'd244, 8'd231}: color_data = 12'h400;
			{9'd244, 8'd232}: color_data = 12'h900;
			{9'd244, 8'd233}: color_data = 12'ha00;
			{9'd244, 8'd234}: color_data = 12'h400;
			{9'd244, 8'd235}: color_data = 12'h310;
			{9'd244, 8'd236}: color_data = 12'hc30;
			{9'd244, 8'd237}: color_data = 12'hc20;
			{9'd244, 8'd238}: color_data = 12'h600;
			{9'd244, 8'd239}: color_data = 12'h000;
			{9'd245, 8'd68}: color_data = 12'h047;
			{9'd245, 8'd69}: color_data = 12'h6df;
			{9'd245, 8'd70}: color_data = 12'hfff;
			{9'd245, 8'd71}: color_data = 12'hcbb;
			{9'd245, 8'd72}: color_data = 12'h323;
			{9'd245, 8'd73}: color_data = 12'h002;
			{9'd245, 8'd74}: color_data = 12'h000;
			{9'd245, 8'd75}: color_data = 12'h012;
			{9'd245, 8'd76}: color_data = 12'h08c;
			{9'd245, 8'd77}: color_data = 12'h034;
			{9'd245, 8'd119}: color_data = 12'h000;
			{9'd245, 8'd120}: color_data = 12'h1ac;
			{9'd245, 8'd121}: color_data = 12'hdff;
			{9'd245, 8'd122}: color_data = 12'hfee;
			{9'd245, 8'd123}: color_data = 12'h666;
			{9'd245, 8'd124}: color_data = 12'h002;
			{9'd245, 8'd125}: color_data = 12'h001;
			{9'd245, 8'd126}: color_data = 12'h000;
			{9'd245, 8'd127}: color_data = 12'h068;
			{9'd245, 8'd128}: color_data = 12'h079;
			{9'd245, 8'd129}: color_data = 12'h000;
			{9'd245, 8'd170}: color_data = 12'h000;
			{9'd245, 8'd171}: color_data = 12'h068;
			{9'd245, 8'd172}: color_data = 12'h8ef;
			{9'd245, 8'd173}: color_data = 12'hfff;
			{9'd245, 8'd174}: color_data = 12'haaa;
			{9'd245, 8'd175}: color_data = 12'h213;
			{9'd245, 8'd176}: color_data = 12'h002;
			{9'd245, 8'd177}: color_data = 12'h000;
			{9'd245, 8'd178}: color_data = 12'h023;
			{9'd245, 8'd179}: color_data = 12'h08c;
			{9'd245, 8'd180}: color_data = 12'h023;
			{9'd245, 8'd222}: color_data = 12'h200;
			{9'd245, 8'd223}: color_data = 12'h900;
			{9'd245, 8'd224}: color_data = 12'ha00;
			{9'd245, 8'd225}: color_data = 12'h800;
			{9'd245, 8'd226}: color_data = 12'h100;
			{9'd245, 8'd227}: color_data = 12'h100;
			{9'd245, 8'd228}: color_data = 12'h310;
			{9'd245, 8'd229}: color_data = 12'h200;
			{9'd245, 8'd230}: color_data = 12'h000;
			{9'd245, 8'd231}: color_data = 12'h500;
			{9'd245, 8'd232}: color_data = 12'ha00;
			{9'd245, 8'd233}: color_data = 12'ha00;
			{9'd245, 8'd234}: color_data = 12'h500;
			{9'd245, 8'd235}: color_data = 12'h000;
			{9'd245, 8'd236}: color_data = 12'h200;
			{9'd245, 8'd237}: color_data = 12'h300;
			{9'd245, 8'd238}: color_data = 12'h100;
			{9'd245, 8'd239}: color_data = 12'h000;
			{9'd246, 8'd68}: color_data = 12'h047;
			{9'd246, 8'd69}: color_data = 12'h6ef;
			{9'd246, 8'd70}: color_data = 12'hddc;
			{9'd246, 8'd71}: color_data = 12'h434;
			{9'd246, 8'd72}: color_data = 12'h003;
			{9'd246, 8'd73}: color_data = 12'h005;
			{9'd246, 8'd74}: color_data = 12'h002;
			{9'd246, 8'd75}: color_data = 12'h012;
			{9'd246, 8'd76}: color_data = 12'h08c;
			{9'd246, 8'd77}: color_data = 12'h034;
			{9'd246, 8'd119}: color_data = 12'h000;
			{9'd246, 8'd120}: color_data = 12'h2ad;
			{9'd246, 8'd121}: color_data = 12'hcff;
			{9'd246, 8'd122}: color_data = 12'h877;
			{9'd246, 8'd123}: color_data = 12'h002;
			{9'd246, 8'd124}: color_data = 12'h004;
			{9'd246, 8'd125}: color_data = 12'h004;
			{9'd246, 8'd126}: color_data = 12'h000;
			{9'd246, 8'd127}: color_data = 12'h068;
			{9'd246, 8'd128}: color_data = 12'h079;
			{9'd246, 8'd129}: color_data = 12'h000;
			{9'd246, 8'd170}: color_data = 12'h000;
			{9'd246, 8'd171}: color_data = 12'h068;
			{9'd246, 8'd172}: color_data = 12'h8ff;
			{9'd246, 8'd173}: color_data = 12'hcbb;
			{9'd246, 8'd174}: color_data = 12'h223;
			{9'd246, 8'd175}: color_data = 12'h003;
			{9'd246, 8'd176}: color_data = 12'h005;
			{9'd246, 8'd177}: color_data = 12'h002;
			{9'd246, 8'd178}: color_data = 12'h023;
			{9'd246, 8'd179}: color_data = 12'h09c;
			{9'd246, 8'd180}: color_data = 12'h023;
			{9'd246, 8'd222}: color_data = 12'h300;
			{9'd246, 8'd223}: color_data = 12'hc20;
			{9'd246, 8'd224}: color_data = 12'ha00;
			{9'd246, 8'd225}: color_data = 12'h800;
			{9'd246, 8'd226}: color_data = 12'h100;
			{9'd246, 8'd227}: color_data = 12'h300;
			{9'd246, 8'd228}: color_data = 12'h500;
			{9'd246, 8'd229}: color_data = 12'h500;
			{9'd246, 8'd230}: color_data = 12'h100;
			{9'd246, 8'd231}: color_data = 12'h710;
			{9'd246, 8'd232}: color_data = 12'hc10;
			{9'd246, 8'd233}: color_data = 12'h900;
			{9'd246, 8'd234}: color_data = 12'h500;
			{9'd246, 8'd235}: color_data = 12'h100;
			{9'd246, 8'd236}: color_data = 12'h500;
			{9'd246, 8'd237}: color_data = 12'h500;
			{9'd246, 8'd238}: color_data = 12'h400;
			{9'd246, 8'd239}: color_data = 12'h000;
			{9'd247, 8'd68}: color_data = 12'h057;
			{9'd247, 8'd69}: color_data = 12'h3bd;
			{9'd247, 8'd70}: color_data = 12'h555;
			{9'd247, 8'd71}: color_data = 12'h002;
			{9'd247, 8'd72}: color_data = 12'h005;
			{9'd247, 8'd73}: color_data = 12'h005;
			{9'd247, 8'd74}: color_data = 12'h004;
			{9'd247, 8'd75}: color_data = 12'h025;
			{9'd247, 8'd76}: color_data = 12'h09c;
			{9'd247, 8'd77}: color_data = 12'h034;
			{9'd247, 8'd119}: color_data = 12'h000;
			{9'd247, 8'd120}: color_data = 12'h1ac;
			{9'd247, 8'd121}: color_data = 12'h699;
			{9'd247, 8'd122}: color_data = 12'h212;
			{9'd247, 8'd123}: color_data = 12'h004;
			{9'd247, 8'd124}: color_data = 12'h005;
			{9'd247, 8'd125}: color_data = 12'h005;
			{9'd247, 8'd126}: color_data = 12'h003;
			{9'd247, 8'd127}: color_data = 12'h06a;
			{9'd247, 8'd128}: color_data = 12'h079;
			{9'd247, 8'd129}: color_data = 12'h000;
			{9'd247, 8'd170}: color_data = 12'h000;
			{9'd247, 8'd171}: color_data = 12'h079;
			{9'd247, 8'd172}: color_data = 12'h4bd;
			{9'd247, 8'd173}: color_data = 12'h444;
			{9'd247, 8'd174}: color_data = 12'h002;
			{9'd247, 8'd175}: color_data = 12'h005;
			{9'd247, 8'd176}: color_data = 12'h005;
			{9'd247, 8'd177}: color_data = 12'h004;
			{9'd247, 8'd178}: color_data = 12'h036;
			{9'd247, 8'd179}: color_data = 12'h09c;
			{9'd247, 8'd180}: color_data = 12'h023;
			{9'd247, 8'd222}: color_data = 12'h410;
			{9'd247, 8'd223}: color_data = 12'hd30;
			{9'd247, 8'd224}: color_data = 12'hb00;
			{9'd247, 8'd225}: color_data = 12'h700;
			{9'd247, 8'd226}: color_data = 12'h200;
			{9'd247, 8'd227}: color_data = 12'h700;
			{9'd247, 8'd228}: color_data = 12'hb00;
			{9'd247, 8'd229}: color_data = 12'h900;
			{9'd247, 8'd230}: color_data = 12'h300;
			{9'd247, 8'd231}: color_data = 12'h820;
			{9'd247, 8'd232}: color_data = 12'hd20;
			{9'd247, 8'd233}: color_data = 12'h900;
			{9'd247, 8'd234}: color_data = 12'h500;
			{9'd247, 8'd235}: color_data = 12'h300;
			{9'd247, 8'd236}: color_data = 12'h900;
			{9'd247, 8'd237}: color_data = 12'hb00;
			{9'd247, 8'd238}: color_data = 12'h800;
			{9'd247, 8'd239}: color_data = 12'h100;
			{9'd248, 8'd68}: color_data = 12'h035;
			{9'd248, 8'd69}: color_data = 12'h047;
			{9'd248, 8'd70}: color_data = 12'h001;
			{9'd248, 8'd71}: color_data = 12'h004;
			{9'd248, 8'd72}: color_data = 12'h004;
			{9'd248, 8'd73}: color_data = 12'h004;
			{9'd248, 8'd74}: color_data = 12'h004;
			{9'd248, 8'd75}: color_data = 12'h015;
			{9'd248, 8'd76}: color_data = 12'h059;
			{9'd248, 8'd77}: color_data = 12'h023;
			{9'd248, 8'd119}: color_data = 12'h000;
			{9'd248, 8'd120}: color_data = 12'h059;
			{9'd248, 8'd121}: color_data = 12'h024;
			{9'd248, 8'd122}: color_data = 12'h004;
			{9'd248, 8'd123}: color_data = 12'h006;
			{9'd248, 8'd124}: color_data = 12'h005;
			{9'd248, 8'd125}: color_data = 12'h005;
			{9'd248, 8'd126}: color_data = 12'h005;
			{9'd248, 8'd127}: color_data = 12'h04a;
			{9'd248, 8'd128}: color_data = 12'h047;
			{9'd248, 8'd129}: color_data = 12'h000;
			{9'd248, 8'd170}: color_data = 12'h000;
			{9'd248, 8'd171}: color_data = 12'h047;
			{9'd248, 8'd172}: color_data = 12'h036;
			{9'd248, 8'd173}: color_data = 12'h001;
			{9'd248, 8'd174}: color_data = 12'h004;
			{9'd248, 8'd175}: color_data = 12'h004;
			{9'd248, 8'd176}: color_data = 12'h004;
			{9'd248, 8'd177}: color_data = 12'h004;
			{9'd248, 8'd178}: color_data = 12'h016;
			{9'd248, 8'd179}: color_data = 12'h059;
			{9'd248, 8'd180}: color_data = 12'h012;
			{9'd248, 8'd222}: color_data = 12'h410;
			{9'd248, 8'd223}: color_data = 12'he40;
			{9'd248, 8'd224}: color_data = 12'hd20;
			{9'd248, 8'd225}: color_data = 12'h800;
			{9'd248, 8'd226}: color_data = 12'h200;
			{9'd248, 8'd227}: color_data = 12'h600;
			{9'd248, 8'd228}: color_data = 12'ha00;
			{9'd248, 8'd229}: color_data = 12'h900;
			{9'd248, 8'd230}: color_data = 12'h300;
			{9'd248, 8'd231}: color_data = 12'h820;
			{9'd248, 8'd232}: color_data = 12'hf30;
			{9'd248, 8'd233}: color_data = 12'hc00;
			{9'd248, 8'd234}: color_data = 12'h500;
			{9'd248, 8'd235}: color_data = 12'h200;
			{9'd248, 8'd236}: color_data = 12'h900;
			{9'd248, 8'd237}: color_data = 12'ha00;
			{9'd248, 8'd238}: color_data = 12'h700;
			{9'd248, 8'd239}: color_data = 12'h100;
			{9'd249, 8'd68}: color_data = 12'h013;
			{9'd249, 8'd69}: color_data = 12'h027;
			{9'd249, 8'd70}: color_data = 12'h016;
			{9'd249, 8'd71}: color_data = 12'h027;
			{9'd249, 8'd72}: color_data = 12'h027;
			{9'd249, 8'd73}: color_data = 12'h017;
			{9'd249, 8'd74}: color_data = 12'h027;
			{9'd249, 8'd75}: color_data = 12'h028;
			{9'd249, 8'd76}: color_data = 12'h027;
			{9'd249, 8'd77}: color_data = 12'h001;
			{9'd249, 8'd119}: color_data = 12'h000;
			{9'd249, 8'd120}: color_data = 12'h003;
			{9'd249, 8'd121}: color_data = 12'h004;
			{9'd249, 8'd122}: color_data = 12'h004;
			{9'd249, 8'd123}: color_data = 12'h004;
			{9'd249, 8'd124}: color_data = 12'h004;
			{9'd249, 8'd125}: color_data = 12'h004;
			{9'd249, 8'd126}: color_data = 12'h004;
			{9'd249, 8'd127}: color_data = 12'h005;
			{9'd249, 8'd128}: color_data = 12'h002;
			{9'd249, 8'd129}: color_data = 12'h000;
			{9'd249, 8'd170}: color_data = 12'h000;
			{9'd249, 8'd171}: color_data = 12'h014;
			{9'd249, 8'd172}: color_data = 12'h027;
			{9'd249, 8'd173}: color_data = 12'h016;
			{9'd249, 8'd174}: color_data = 12'h027;
			{9'd249, 8'd175}: color_data = 12'h027;
			{9'd249, 8'd176}: color_data = 12'h017;
			{9'd249, 8'd177}: color_data = 12'h027;
			{9'd249, 8'd178}: color_data = 12'h028;
			{9'd249, 8'd179}: color_data = 12'h026;
			{9'd249, 8'd180}: color_data = 12'h001;
			{9'd249, 8'd222}: color_data = 12'h300;
			{9'd249, 8'd223}: color_data = 12'hc30;
			{9'd249, 8'd224}: color_data = 12'hc30;
			{9'd249, 8'd225}: color_data = 12'h600;
			{9'd249, 8'd226}: color_data = 12'h100;
			{9'd249, 8'd227}: color_data = 12'h600;
			{9'd249, 8'd228}: color_data = 12'ha00;
			{9'd249, 8'd229}: color_data = 12'h900;
			{9'd249, 8'd230}: color_data = 12'h300;
			{9'd249, 8'd231}: color_data = 12'h620;
			{9'd249, 8'd232}: color_data = 12'hd40;
			{9'd249, 8'd233}: color_data = 12'ha20;
			{9'd249, 8'd234}: color_data = 12'h300;
			{9'd249, 8'd235}: color_data = 12'h200;
			{9'd249, 8'd236}: color_data = 12'h900;
			{9'd249, 8'd237}: color_data = 12'ha00;
			{9'd249, 8'd238}: color_data = 12'h700;
			{9'd249, 8'd239}: color_data = 12'h100;
			{9'd250, 8'd68}: color_data = 12'h035;
			{9'd250, 8'd69}: color_data = 12'h09e;
			{9'd250, 8'd70}: color_data = 12'h09e;
			{9'd250, 8'd71}: color_data = 12'h09e;
			{9'd250, 8'd72}: color_data = 12'h09e;
			{9'd250, 8'd73}: color_data = 12'h09e;
			{9'd250, 8'd74}: color_data = 12'h09e;
			{9'd250, 8'd75}: color_data = 12'h09e;
			{9'd250, 8'd76}: color_data = 12'h08c;
			{9'd250, 8'd77}: color_data = 12'h023;
			{9'd250, 8'd120}: color_data = 12'h000;
			{9'd250, 8'd121}: color_data = 12'h001;
			{9'd250, 8'd122}: color_data = 12'h001;
			{9'd250, 8'd123}: color_data = 12'h000;
			{9'd250, 8'd124}: color_data = 12'h000;
			{9'd250, 8'd125}: color_data = 12'h000;
			{9'd250, 8'd126}: color_data = 12'h000;
			{9'd250, 8'd127}: color_data = 12'h000;
			{9'd250, 8'd128}: color_data = 12'h000;
			{9'd250, 8'd170}: color_data = 12'h000;
			{9'd250, 8'd171}: color_data = 12'h057;
			{9'd250, 8'd172}: color_data = 12'h0ae;
			{9'd250, 8'd173}: color_data = 12'h09e;
			{9'd250, 8'd174}: color_data = 12'h09e;
			{9'd250, 8'd175}: color_data = 12'h09e;
			{9'd250, 8'd176}: color_data = 12'h09e;
			{9'd250, 8'd177}: color_data = 12'h09e;
			{9'd250, 8'd178}: color_data = 12'h09e;
			{9'd250, 8'd179}: color_data = 12'h07b;
			{9'd250, 8'd180}: color_data = 12'h012;
			{9'd250, 8'd222}: color_data = 12'h000;
			{9'd250, 8'd223}: color_data = 12'h200;
			{9'd250, 8'd224}: color_data = 12'h300;
			{9'd250, 8'd225}: color_data = 12'h100;
			{9'd250, 8'd226}: color_data = 12'h000;
			{9'd250, 8'd227}: color_data = 12'h700;
			{9'd250, 8'd228}: color_data = 12'ha00;
			{9'd250, 8'd229}: color_data = 12'h900;
			{9'd250, 8'd230}: color_data = 12'h300;
			{9'd250, 8'd231}: color_data = 12'h100;
			{9'd250, 8'd232}: color_data = 12'h310;
			{9'd250, 8'd233}: color_data = 12'h200;
			{9'd250, 8'd234}: color_data = 12'h000;
			{9'd250, 8'd235}: color_data = 12'h300;
			{9'd250, 8'd236}: color_data = 12'h900;
			{9'd250, 8'd237}: color_data = 12'ha00;
			{9'd250, 8'd238}: color_data = 12'h700;
			{9'd250, 8'd239}: color_data = 12'h100;
			{9'd251, 8'd68}: color_data = 12'h057;
			{9'd251, 8'd69}: color_data = 12'h4ef;
			{9'd251, 8'd70}: color_data = 12'h7ef;
			{9'd251, 8'd71}: color_data = 12'h0cf;
			{9'd251, 8'd72}: color_data = 12'h0cf;
			{9'd251, 8'd73}: color_data = 12'h0df;
			{9'd251, 8'd74}: color_data = 12'h0bd;
			{9'd251, 8'd75}: color_data = 12'h068;
			{9'd251, 8'd76}: color_data = 12'h09c;
			{9'd251, 8'd77}: color_data = 12'h034;
			{9'd251, 8'd170}: color_data = 12'h000;
			{9'd251, 8'd171}: color_data = 12'h069;
			{9'd251, 8'd172}: color_data = 12'h6ef;
			{9'd251, 8'd173}: color_data = 12'h6ef;
			{9'd251, 8'd174}: color_data = 12'h0cf;
			{9'd251, 8'd175}: color_data = 12'h0cf;
			{9'd251, 8'd176}: color_data = 12'h0df;
			{9'd251, 8'd177}: color_data = 12'h0ac;
			{9'd251, 8'd178}: color_data = 12'h079;
			{9'd251, 8'd179}: color_data = 12'h09c;
			{9'd251, 8'd180}: color_data = 12'h023;
			{9'd251, 8'd222}: color_data = 12'h100;
			{9'd251, 8'd223}: color_data = 12'h500;
			{9'd251, 8'd224}: color_data = 12'h600;
			{9'd251, 8'd225}: color_data = 12'h400;
			{9'd251, 8'd226}: color_data = 12'h100;
			{9'd251, 8'd227}: color_data = 12'ha20;
			{9'd251, 8'd228}: color_data = 12'hb10;
			{9'd251, 8'd229}: color_data = 12'h900;
			{9'd251, 8'd230}: color_data = 12'h300;
			{9'd251, 8'd231}: color_data = 12'h200;
			{9'd251, 8'd232}: color_data = 12'h500;
			{9'd251, 8'd233}: color_data = 12'h500;
			{9'd251, 8'd234}: color_data = 12'h200;
			{9'd251, 8'd235}: color_data = 12'h410;
			{9'd251, 8'd236}: color_data = 12'hc20;
			{9'd251, 8'd237}: color_data = 12'ha00;
			{9'd251, 8'd238}: color_data = 12'h700;
			{9'd251, 8'd239}: color_data = 12'h100;
			{9'd252, 8'd68}: color_data = 12'h047;
			{9'd252, 8'd69}: color_data = 12'h6df;
			{9'd252, 8'd70}: color_data = 12'heff;
			{9'd252, 8'd71}: color_data = 12'h6df;
			{9'd252, 8'd72}: color_data = 12'h0bf;
			{9'd252, 8'd73}: color_data = 12'h0bf;
			{9'd252, 8'd74}: color_data = 12'h056;
			{9'd252, 8'd75}: color_data = 12'h012;
			{9'd252, 8'd76}: color_data = 12'h08b;
			{9'd252, 8'd77}: color_data = 12'h034;
			{9'd252, 8'd170}: color_data = 12'h000;
			{9'd252, 8'd171}: color_data = 12'h068;
			{9'd252, 8'd172}: color_data = 12'h8ef;
			{9'd252, 8'd173}: color_data = 12'hdff;
			{9'd252, 8'd174}: color_data = 12'h4cf;
			{9'd252, 8'd175}: color_data = 12'h0cf;
			{9'd252, 8'd176}: color_data = 12'h0ae;
			{9'd252, 8'd177}: color_data = 12'h035;
			{9'd252, 8'd178}: color_data = 12'h023;
			{9'd252, 8'd179}: color_data = 12'h08c;
			{9'd252, 8'd180}: color_data = 12'h023;
			{9'd252, 8'd222}: color_data = 12'h200;
			{9'd252, 8'd223}: color_data = 12'h900;
			{9'd252, 8'd224}: color_data = 12'hb00;
			{9'd252, 8'd225}: color_data = 12'h800;
			{9'd252, 8'd226}: color_data = 12'h200;
			{9'd252, 8'd227}: color_data = 12'hb30;
			{9'd252, 8'd228}: color_data = 12'hc10;
			{9'd252, 8'd229}: color_data = 12'h800;
			{9'd252, 8'd230}: color_data = 12'h300;
			{9'd252, 8'd231}: color_data = 12'h500;
			{9'd252, 8'd232}: color_data = 12'ha00;
			{9'd252, 8'd233}: color_data = 12'ha00;
			{9'd252, 8'd234}: color_data = 12'h500;
			{9'd252, 8'd235}: color_data = 12'h510;
			{9'd252, 8'd236}: color_data = 12'hd30;
			{9'd252, 8'd237}: color_data = 12'ha00;
			{9'd252, 8'd238}: color_data = 12'h700;
			{9'd252, 8'd239}: color_data = 12'h100;
			{9'd253, 8'd68}: color_data = 12'h047;
			{9'd253, 8'd69}: color_data = 12'h6df;
			{9'd253, 8'd70}: color_data = 12'hfff;
			{9'd253, 8'd71}: color_data = 12'hdff;
			{9'd253, 8'd72}: color_data = 12'h5df;
			{9'd253, 8'd73}: color_data = 12'h068;
			{9'd253, 8'd74}: color_data = 12'h000;
			{9'd253, 8'd75}: color_data = 12'h012;
			{9'd253, 8'd76}: color_data = 12'h08c;
			{9'd253, 8'd77}: color_data = 12'h034;
			{9'd253, 8'd170}: color_data = 12'h000;
			{9'd253, 8'd171}: color_data = 12'h068;
			{9'd253, 8'd172}: color_data = 12'h8ef;
			{9'd253, 8'd173}: color_data = 12'hfff;
			{9'd253, 8'd174}: color_data = 12'hcff;
			{9'd253, 8'd175}: color_data = 12'h4ce;
			{9'd253, 8'd176}: color_data = 12'h057;
			{9'd253, 8'd177}: color_data = 12'h000;
			{9'd253, 8'd178}: color_data = 12'h023;
			{9'd253, 8'd179}: color_data = 12'h08c;
			{9'd253, 8'd180}: color_data = 12'h023;
			{9'd253, 8'd222}: color_data = 12'h200;
			{9'd253, 8'd223}: color_data = 12'h900;
			{9'd253, 8'd224}: color_data = 12'ha00;
			{9'd253, 8'd225}: color_data = 12'h700;
			{9'd253, 8'd226}: color_data = 12'h200;
			{9'd253, 8'd227}: color_data = 12'hb30;
			{9'd253, 8'd228}: color_data = 12'he20;
			{9'd253, 8'd229}: color_data = 12'ha00;
			{9'd253, 8'd230}: color_data = 12'h300;
			{9'd253, 8'd231}: color_data = 12'h400;
			{9'd253, 8'd232}: color_data = 12'ha00;
			{9'd253, 8'd233}: color_data = 12'ha00;
			{9'd253, 8'd234}: color_data = 12'h400;
			{9'd253, 8'd235}: color_data = 12'h510;
			{9'd253, 8'd236}: color_data = 12'hf40;
			{9'd253, 8'd237}: color_data = 12'hd10;
			{9'd253, 8'd238}: color_data = 12'h800;
			{9'd253, 8'd239}: color_data = 12'h100;
			{9'd254, 8'd68}: color_data = 12'h047;
			{9'd254, 8'd69}: color_data = 12'h6df;
			{9'd254, 8'd70}: color_data = 12'hfff;
			{9'd254, 8'd71}: color_data = 12'hfff;
			{9'd254, 8'd72}: color_data = 12'h9aa;
			{9'd254, 8'd73}: color_data = 12'h011;
			{9'd254, 8'd75}: color_data = 12'h012;
			{9'd254, 8'd76}: color_data = 12'h08c;
			{9'd254, 8'd77}: color_data = 12'h034;
			{9'd254, 8'd170}: color_data = 12'h000;
			{9'd254, 8'd171}: color_data = 12'h068;
			{9'd254, 8'd172}: color_data = 12'h7ef;
			{9'd254, 8'd173}: color_data = 12'hfff;
			{9'd254, 8'd174}: color_data = 12'hfff;
			{9'd254, 8'd175}: color_data = 12'h899;
			{9'd254, 8'd176}: color_data = 12'h001;
			{9'd254, 8'd178}: color_data = 12'h024;
			{9'd254, 8'd179}: color_data = 12'h08c;
			{9'd254, 8'd180}: color_data = 12'h023;
			{9'd254, 8'd222}: color_data = 12'h200;
			{9'd254, 8'd223}: color_data = 12'h800;
			{9'd254, 8'd224}: color_data = 12'ha00;
			{9'd254, 8'd225}: color_data = 12'h800;
			{9'd254, 8'd226}: color_data = 12'h200;
			{9'd254, 8'd227}: color_data = 12'h920;
			{9'd254, 8'd228}: color_data = 12'hd30;
			{9'd254, 8'd229}: color_data = 12'h910;
			{9'd254, 8'd230}: color_data = 12'h200;
			{9'd254, 8'd231}: color_data = 12'h400;
			{9'd254, 8'd232}: color_data = 12'h900;
			{9'd254, 8'd233}: color_data = 12'ha00;
			{9'd254, 8'd234}: color_data = 12'h400;
			{9'd254, 8'd235}: color_data = 12'h310;
			{9'd254, 8'd236}: color_data = 12'hc30;
			{9'd254, 8'd237}: color_data = 12'hc20;
			{9'd254, 8'd238}: color_data = 12'h600;
			{9'd254, 8'd239}: color_data = 12'h000;
			{9'd255, 8'd68}: color_data = 12'h047;
			{9'd255, 8'd69}: color_data = 12'h6df;
			{9'd255, 8'd70}: color_data = 12'hfff;
			{9'd255, 8'd71}: color_data = 12'hcbb;
			{9'd255, 8'd72}: color_data = 12'h323;
			{9'd255, 8'd73}: color_data = 12'h002;
			{9'd255, 8'd74}: color_data = 12'h000;
			{9'd255, 8'd75}: color_data = 12'h012;
			{9'd255, 8'd76}: color_data = 12'h08c;
			{9'd255, 8'd77}: color_data = 12'h034;
			{9'd255, 8'd170}: color_data = 12'h000;
			{9'd255, 8'd171}: color_data = 12'h068;
			{9'd255, 8'd172}: color_data = 12'h8ef;
			{9'd255, 8'd173}: color_data = 12'hfff;
			{9'd255, 8'd174}: color_data = 12'haa9;
			{9'd255, 8'd175}: color_data = 12'h212;
			{9'd255, 8'd176}: color_data = 12'h002;
			{9'd255, 8'd177}: color_data = 12'h000;
			{9'd255, 8'd178}: color_data = 12'h023;
			{9'd255, 8'd179}: color_data = 12'h08c;
			{9'd255, 8'd180}: color_data = 12'h023;
			{9'd255, 8'd222}: color_data = 12'h200;
			{9'd255, 8'd223}: color_data = 12'h900;
			{9'd255, 8'd224}: color_data = 12'ha00;
			{9'd255, 8'd225}: color_data = 12'h800;
			{9'd255, 8'd226}: color_data = 12'h100;
			{9'd255, 8'd227}: color_data = 12'h100;
			{9'd255, 8'd228}: color_data = 12'h310;
			{9'd255, 8'd229}: color_data = 12'h200;
			{9'd255, 8'd230}: color_data = 12'h000;
			{9'd255, 8'd231}: color_data = 12'h500;
			{9'd255, 8'd232}: color_data = 12'ha00;
			{9'd255, 8'd233}: color_data = 12'ha00;
			{9'd255, 8'd234}: color_data = 12'h500;
			{9'd255, 8'd235}: color_data = 12'h000;
			{9'd255, 8'd236}: color_data = 12'h200;
			{9'd255, 8'd237}: color_data = 12'h300;
			{9'd255, 8'd238}: color_data = 12'h100;
			{9'd255, 8'd239}: color_data = 12'h000;
			{9'd256, 8'd68}: color_data = 12'h047;
			{9'd256, 8'd69}: color_data = 12'h6ef;
			{9'd256, 8'd70}: color_data = 12'hdcc;
			{9'd256, 8'd71}: color_data = 12'h434;
			{9'd256, 8'd72}: color_data = 12'h003;
			{9'd256, 8'd73}: color_data = 12'h005;
			{9'd256, 8'd74}: color_data = 12'h002;
			{9'd256, 8'd75}: color_data = 12'h012;
			{9'd256, 8'd76}: color_data = 12'h08c;
			{9'd256, 8'd77}: color_data = 12'h034;
			{9'd256, 8'd170}: color_data = 12'h000;
			{9'd256, 8'd171}: color_data = 12'h068;
			{9'd256, 8'd172}: color_data = 12'h8ff;
			{9'd256, 8'd173}: color_data = 12'hcbb;
			{9'd256, 8'd174}: color_data = 12'h323;
			{9'd256, 8'd175}: color_data = 12'h003;
			{9'd256, 8'd176}: color_data = 12'h005;
			{9'd256, 8'd177}: color_data = 12'h002;
			{9'd256, 8'd178}: color_data = 12'h023;
			{9'd256, 8'd179}: color_data = 12'h09c;
			{9'd256, 8'd180}: color_data = 12'h023;
			{9'd256, 8'd222}: color_data = 12'h300;
			{9'd256, 8'd223}: color_data = 12'hc20;
			{9'd256, 8'd224}: color_data = 12'ha00;
			{9'd256, 8'd225}: color_data = 12'h800;
			{9'd256, 8'd226}: color_data = 12'h100;
			{9'd256, 8'd227}: color_data = 12'h300;
			{9'd256, 8'd228}: color_data = 12'h500;
			{9'd256, 8'd229}: color_data = 12'h500;
			{9'd256, 8'd230}: color_data = 12'h100;
			{9'd256, 8'd231}: color_data = 12'h710;
			{9'd256, 8'd232}: color_data = 12'hc10;
			{9'd256, 8'd233}: color_data = 12'h900;
			{9'd256, 8'd234}: color_data = 12'h500;
			{9'd256, 8'd235}: color_data = 12'h100;
			{9'd256, 8'd236}: color_data = 12'h500;
			{9'd256, 8'd237}: color_data = 12'h600;
			{9'd256, 8'd238}: color_data = 12'h400;
			{9'd256, 8'd239}: color_data = 12'h000;
			{9'd257, 8'd68}: color_data = 12'h057;
			{9'd257, 8'd69}: color_data = 12'h3bd;
			{9'd257, 8'd70}: color_data = 12'h555;
			{9'd257, 8'd71}: color_data = 12'h002;
			{9'd257, 8'd72}: color_data = 12'h005;
			{9'd257, 8'd73}: color_data = 12'h005;
			{9'd257, 8'd74}: color_data = 12'h004;
			{9'd257, 8'd75}: color_data = 12'h025;
			{9'd257, 8'd76}: color_data = 12'h09c;
			{9'd257, 8'd77}: color_data = 12'h034;
			{9'd257, 8'd170}: color_data = 12'h000;
			{9'd257, 8'd171}: color_data = 12'h079;
			{9'd257, 8'd172}: color_data = 12'h4bd;
			{9'd257, 8'd173}: color_data = 12'h444;
			{9'd257, 8'd174}: color_data = 12'h002;
			{9'd257, 8'd175}: color_data = 12'h005;
			{9'd257, 8'd176}: color_data = 12'h005;
			{9'd257, 8'd177}: color_data = 12'h004;
			{9'd257, 8'd178}: color_data = 12'h036;
			{9'd257, 8'd179}: color_data = 12'h09c;
			{9'd257, 8'd180}: color_data = 12'h023;
			{9'd257, 8'd222}: color_data = 12'h410;
			{9'd257, 8'd223}: color_data = 12'hd30;
			{9'd257, 8'd224}: color_data = 12'hb00;
			{9'd257, 8'd225}: color_data = 12'h700;
			{9'd257, 8'd226}: color_data = 12'h200;
			{9'd257, 8'd227}: color_data = 12'h700;
			{9'd257, 8'd228}: color_data = 12'hb00;
			{9'd257, 8'd229}: color_data = 12'ha00;
			{9'd257, 8'd230}: color_data = 12'h300;
			{9'd257, 8'd231}: color_data = 12'h820;
			{9'd257, 8'd232}: color_data = 12'hd20;
			{9'd257, 8'd233}: color_data = 12'h900;
			{9'd257, 8'd234}: color_data = 12'h500;
			{9'd257, 8'd235}: color_data = 12'h300;
			{9'd257, 8'd236}: color_data = 12'h900;
			{9'd257, 8'd237}: color_data = 12'hb00;
			{9'd257, 8'd238}: color_data = 12'h800;
			{9'd257, 8'd239}: color_data = 12'h100;
			{9'd258, 8'd68}: color_data = 12'h035;
			{9'd258, 8'd69}: color_data = 12'h047;
			{9'd258, 8'd70}: color_data = 12'h001;
			{9'd258, 8'd71}: color_data = 12'h004;
			{9'd258, 8'd72}: color_data = 12'h004;
			{9'd258, 8'd73}: color_data = 12'h004;
			{9'd258, 8'd74}: color_data = 12'h004;
			{9'd258, 8'd75}: color_data = 12'h015;
			{9'd258, 8'd76}: color_data = 12'h059;
			{9'd258, 8'd77}: color_data = 12'h023;
			{9'd258, 8'd170}: color_data = 12'h000;
			{9'd258, 8'd171}: color_data = 12'h047;
			{9'd258, 8'd172}: color_data = 12'h036;
			{9'd258, 8'd173}: color_data = 12'h001;
			{9'd258, 8'd174}: color_data = 12'h004;
			{9'd258, 8'd175}: color_data = 12'h004;
			{9'd258, 8'd176}: color_data = 12'h004;
			{9'd258, 8'd177}: color_data = 12'h004;
			{9'd258, 8'd178}: color_data = 12'h016;
			{9'd258, 8'd179}: color_data = 12'h059;
			{9'd258, 8'd180}: color_data = 12'h012;
			{9'd258, 8'd222}: color_data = 12'h410;
			{9'd258, 8'd223}: color_data = 12'he40;
			{9'd258, 8'd224}: color_data = 12'hd20;
			{9'd258, 8'd225}: color_data = 12'h800;
			{9'd258, 8'd226}: color_data = 12'h200;
			{9'd258, 8'd227}: color_data = 12'h600;
			{9'd258, 8'd228}: color_data = 12'ha00;
			{9'd258, 8'd229}: color_data = 12'h900;
			{9'd258, 8'd230}: color_data = 12'h300;
			{9'd258, 8'd231}: color_data = 12'h820;
			{9'd258, 8'd232}: color_data = 12'hf30;
			{9'd258, 8'd233}: color_data = 12'hc00;
			{9'd258, 8'd234}: color_data = 12'h500;
			{9'd258, 8'd235}: color_data = 12'h200;
			{9'd258, 8'd236}: color_data = 12'h900;
			{9'd258, 8'd237}: color_data = 12'ha00;
			{9'd258, 8'd238}: color_data = 12'h700;
			{9'd258, 8'd239}: color_data = 12'h100;
			{9'd259, 8'd68}: color_data = 12'h013;
			{9'd259, 8'd69}: color_data = 12'h027;
			{9'd259, 8'd70}: color_data = 12'h016;
			{9'd259, 8'd71}: color_data = 12'h027;
			{9'd259, 8'd72}: color_data = 12'h027;
			{9'd259, 8'd73}: color_data = 12'h027;
			{9'd259, 8'd74}: color_data = 12'h027;
			{9'd259, 8'd75}: color_data = 12'h028;
			{9'd259, 8'd76}: color_data = 12'h027;
			{9'd259, 8'd77}: color_data = 12'h001;
			{9'd259, 8'd170}: color_data = 12'h000;
			{9'd259, 8'd171}: color_data = 12'h014;
			{9'd259, 8'd172}: color_data = 12'h027;
			{9'd259, 8'd173}: color_data = 12'h016;
			{9'd259, 8'd174}: color_data = 12'h027;
			{9'd259, 8'd175}: color_data = 12'h027;
			{9'd259, 8'd176}: color_data = 12'h026;
			{9'd259, 8'd177}: color_data = 12'h027;
			{9'd259, 8'd178}: color_data = 12'h028;
			{9'd259, 8'd179}: color_data = 12'h026;
			{9'd259, 8'd180}: color_data = 12'h001;
			{9'd259, 8'd222}: color_data = 12'h300;
			{9'd259, 8'd223}: color_data = 12'hc30;
			{9'd259, 8'd224}: color_data = 12'hc30;
			{9'd259, 8'd225}: color_data = 12'h600;
			{9'd259, 8'd226}: color_data = 12'h100;
			{9'd259, 8'd227}: color_data = 12'h600;
			{9'd259, 8'd228}: color_data = 12'ha00;
			{9'd259, 8'd229}: color_data = 12'h900;
			{9'd259, 8'd230}: color_data = 12'h300;
			{9'd259, 8'd231}: color_data = 12'h620;
			{9'd259, 8'd232}: color_data = 12'hd40;
			{9'd259, 8'd233}: color_data = 12'ha20;
			{9'd259, 8'd234}: color_data = 12'h300;
			{9'd259, 8'd235}: color_data = 12'h200;
			{9'd259, 8'd236}: color_data = 12'h900;
			{9'd259, 8'd237}: color_data = 12'ha00;
			{9'd259, 8'd238}: color_data = 12'h700;
			{9'd259, 8'd239}: color_data = 12'h100;
			{9'd260, 8'd68}: color_data = 12'h036;
			{9'd260, 8'd69}: color_data = 12'h09e;
			{9'd260, 8'd70}: color_data = 12'h09e;
			{9'd260, 8'd71}: color_data = 12'h09e;
			{9'd260, 8'd72}: color_data = 12'h09e;
			{9'd260, 8'd73}: color_data = 12'h09e;
			{9'd260, 8'd74}: color_data = 12'h09e;
			{9'd260, 8'd75}: color_data = 12'h09e;
			{9'd260, 8'd76}: color_data = 12'h08c;
			{9'd260, 8'd77}: color_data = 12'h023;
			{9'd260, 8'd170}: color_data = 12'h000;
			{9'd260, 8'd171}: color_data = 12'h057;
			{9'd260, 8'd172}: color_data = 12'h0ae;
			{9'd260, 8'd173}: color_data = 12'h09e;
			{9'd260, 8'd174}: color_data = 12'h09e;
			{9'd260, 8'd175}: color_data = 12'h09e;
			{9'd260, 8'd176}: color_data = 12'h09e;
			{9'd260, 8'd177}: color_data = 12'h09e;
			{9'd260, 8'd178}: color_data = 12'h09e;
			{9'd260, 8'd179}: color_data = 12'h07b;
			{9'd260, 8'd180}: color_data = 12'h012;
			{9'd260, 8'd222}: color_data = 12'h000;
			{9'd260, 8'd223}: color_data = 12'h200;
			{9'd260, 8'd224}: color_data = 12'h300;
			{9'd260, 8'd225}: color_data = 12'h100;
			{9'd260, 8'd226}: color_data = 12'h000;
			{9'd260, 8'd227}: color_data = 12'h700;
			{9'd260, 8'd228}: color_data = 12'ha00;
			{9'd260, 8'd229}: color_data = 12'h900;
			{9'd260, 8'd230}: color_data = 12'h300;
			{9'd260, 8'd231}: color_data = 12'h100;
			{9'd260, 8'd232}: color_data = 12'h310;
			{9'd260, 8'd233}: color_data = 12'h200;
			{9'd260, 8'd234}: color_data = 12'h000;
			{9'd260, 8'd235}: color_data = 12'h300;
			{9'd260, 8'd236}: color_data = 12'h900;
			{9'd260, 8'd237}: color_data = 12'ha00;
			{9'd260, 8'd238}: color_data = 12'h700;
			{9'd260, 8'd239}: color_data = 12'h100;
			{9'd261, 8'd68}: color_data = 12'h057;
			{9'd261, 8'd69}: color_data = 12'h4ef;
			{9'd261, 8'd70}: color_data = 12'h7ef;
			{9'd261, 8'd71}: color_data = 12'h0cf;
			{9'd261, 8'd72}: color_data = 12'h0cf;
			{9'd261, 8'd73}: color_data = 12'h0df;
			{9'd261, 8'd74}: color_data = 12'h0bd;
			{9'd261, 8'd75}: color_data = 12'h068;
			{9'd261, 8'd76}: color_data = 12'h09c;
			{9'd261, 8'd77}: color_data = 12'h034;
			{9'd261, 8'd170}: color_data = 12'h000;
			{9'd261, 8'd171}: color_data = 12'h069;
			{9'd261, 8'd172}: color_data = 12'h6ef;
			{9'd261, 8'd173}: color_data = 12'h6ef;
			{9'd261, 8'd174}: color_data = 12'h0cf;
			{9'd261, 8'd175}: color_data = 12'h0cf;
			{9'd261, 8'd176}: color_data = 12'h0df;
			{9'd261, 8'd177}: color_data = 12'h0ac;
			{9'd261, 8'd178}: color_data = 12'h079;
			{9'd261, 8'd179}: color_data = 12'h09c;
			{9'd261, 8'd180}: color_data = 12'h023;
			{9'd261, 8'd222}: color_data = 12'h100;
			{9'd261, 8'd223}: color_data = 12'h500;
			{9'd261, 8'd224}: color_data = 12'h600;
			{9'd261, 8'd225}: color_data = 12'h400;
			{9'd261, 8'd226}: color_data = 12'h200;
			{9'd261, 8'd227}: color_data = 12'ha20;
			{9'd261, 8'd228}: color_data = 12'hb10;
			{9'd261, 8'd229}: color_data = 12'h900;
			{9'd261, 8'd230}: color_data = 12'h300;
			{9'd261, 8'd231}: color_data = 12'h200;
			{9'd261, 8'd232}: color_data = 12'h500;
			{9'd261, 8'd233}: color_data = 12'h500;
			{9'd261, 8'd234}: color_data = 12'h200;
			{9'd261, 8'd235}: color_data = 12'h410;
			{9'd261, 8'd236}: color_data = 12'hc20;
			{9'd261, 8'd237}: color_data = 12'ha00;
			{9'd261, 8'd238}: color_data = 12'h700;
			{9'd261, 8'd239}: color_data = 12'h100;
			{9'd262, 8'd68}: color_data = 12'h047;
			{9'd262, 8'd69}: color_data = 12'h6df;
			{9'd262, 8'd70}: color_data = 12'heff;
			{9'd262, 8'd71}: color_data = 12'h6df;
			{9'd262, 8'd72}: color_data = 12'h0bf;
			{9'd262, 8'd73}: color_data = 12'h0be;
			{9'd262, 8'd74}: color_data = 12'h056;
			{9'd262, 8'd75}: color_data = 12'h012;
			{9'd262, 8'd76}: color_data = 12'h08b;
			{9'd262, 8'd77}: color_data = 12'h034;
			{9'd262, 8'd170}: color_data = 12'h000;
			{9'd262, 8'd171}: color_data = 12'h068;
			{9'd262, 8'd172}: color_data = 12'h8ef;
			{9'd262, 8'd173}: color_data = 12'hdff;
			{9'd262, 8'd174}: color_data = 12'h4cf;
			{9'd262, 8'd175}: color_data = 12'h0cf;
			{9'd262, 8'd176}: color_data = 12'h0ae;
			{9'd262, 8'd177}: color_data = 12'h035;
			{9'd262, 8'd178}: color_data = 12'h023;
			{9'd262, 8'd179}: color_data = 12'h08c;
			{9'd262, 8'd180}: color_data = 12'h023;
			{9'd262, 8'd222}: color_data = 12'h200;
			{9'd262, 8'd223}: color_data = 12'h900;
			{9'd262, 8'd224}: color_data = 12'hb00;
			{9'd262, 8'd225}: color_data = 12'h800;
			{9'd262, 8'd226}: color_data = 12'h200;
			{9'd262, 8'd227}: color_data = 12'hb30;
			{9'd262, 8'd228}: color_data = 12'hc10;
			{9'd262, 8'd229}: color_data = 12'h800;
			{9'd262, 8'd230}: color_data = 12'h300;
			{9'd262, 8'd231}: color_data = 12'h400;
			{9'd262, 8'd232}: color_data = 12'ha00;
			{9'd262, 8'd233}: color_data = 12'ha00;
			{9'd262, 8'd234}: color_data = 12'h500;
			{9'd262, 8'd235}: color_data = 12'h510;
			{9'd262, 8'd236}: color_data = 12'hd30;
			{9'd262, 8'd237}: color_data = 12'ha00;
			{9'd262, 8'd238}: color_data = 12'h700;
			{9'd262, 8'd239}: color_data = 12'h100;
			{9'd263, 8'd68}: color_data = 12'h047;
			{9'd263, 8'd69}: color_data = 12'h6df;
			{9'd263, 8'd70}: color_data = 12'hfff;
			{9'd263, 8'd71}: color_data = 12'hdff;
			{9'd263, 8'd72}: color_data = 12'h5df;
			{9'd263, 8'd73}: color_data = 12'h068;
			{9'd263, 8'd74}: color_data = 12'h000;
			{9'd263, 8'd75}: color_data = 12'h012;
			{9'd263, 8'd76}: color_data = 12'h08c;
			{9'd263, 8'd77}: color_data = 12'h034;
			{9'd263, 8'd170}: color_data = 12'h000;
			{9'd263, 8'd171}: color_data = 12'h068;
			{9'd263, 8'd172}: color_data = 12'h8ef;
			{9'd263, 8'd173}: color_data = 12'hfff;
			{9'd263, 8'd174}: color_data = 12'hcff;
			{9'd263, 8'd175}: color_data = 12'h4ce;
			{9'd263, 8'd176}: color_data = 12'h057;
			{9'd263, 8'd177}: color_data = 12'h000;
			{9'd263, 8'd178}: color_data = 12'h023;
			{9'd263, 8'd179}: color_data = 12'h08c;
			{9'd263, 8'd180}: color_data = 12'h023;
			{9'd263, 8'd222}: color_data = 12'h200;
			{9'd263, 8'd223}: color_data = 12'h900;
			{9'd263, 8'd224}: color_data = 12'ha00;
			{9'd263, 8'd225}: color_data = 12'h700;
			{9'd263, 8'd226}: color_data = 12'h200;
			{9'd263, 8'd227}: color_data = 12'hb30;
			{9'd263, 8'd228}: color_data = 12'he20;
			{9'd263, 8'd229}: color_data = 12'ha00;
			{9'd263, 8'd230}: color_data = 12'h300;
			{9'd263, 8'd231}: color_data = 12'h400;
			{9'd263, 8'd232}: color_data = 12'ha00;
			{9'd263, 8'd233}: color_data = 12'ha00;
			{9'd263, 8'd234}: color_data = 12'h400;
			{9'd263, 8'd235}: color_data = 12'h510;
			{9'd263, 8'd236}: color_data = 12'hf40;
			{9'd263, 8'd237}: color_data = 12'hd10;
			{9'd263, 8'd238}: color_data = 12'h800;
			{9'd263, 8'd239}: color_data = 12'h100;
			{9'd264, 8'd68}: color_data = 12'h047;
			{9'd264, 8'd69}: color_data = 12'h6df;
			{9'd264, 8'd70}: color_data = 12'hfff;
			{9'd264, 8'd71}: color_data = 12'hfff;
			{9'd264, 8'd72}: color_data = 12'h9aa;
			{9'd264, 8'd73}: color_data = 12'h011;
			{9'd264, 8'd75}: color_data = 12'h012;
			{9'd264, 8'd76}: color_data = 12'h08c;
			{9'd264, 8'd77}: color_data = 12'h034;
			{9'd264, 8'd170}: color_data = 12'h000;
			{9'd264, 8'd171}: color_data = 12'h068;
			{9'd264, 8'd172}: color_data = 12'h7ef;
			{9'd264, 8'd173}: color_data = 12'hfff;
			{9'd264, 8'd174}: color_data = 12'hfff;
			{9'd264, 8'd175}: color_data = 12'h899;
			{9'd264, 8'd176}: color_data = 12'h001;
			{9'd264, 8'd178}: color_data = 12'h024;
			{9'd264, 8'd179}: color_data = 12'h08c;
			{9'd264, 8'd180}: color_data = 12'h023;
			{9'd264, 8'd222}: color_data = 12'h200;
			{9'd264, 8'd223}: color_data = 12'h800;
			{9'd264, 8'd224}: color_data = 12'ha00;
			{9'd264, 8'd225}: color_data = 12'h700;
			{9'd264, 8'd226}: color_data = 12'h200;
			{9'd264, 8'd227}: color_data = 12'h920;
			{9'd264, 8'd228}: color_data = 12'hd30;
			{9'd264, 8'd229}: color_data = 12'h910;
			{9'd264, 8'd230}: color_data = 12'h200;
			{9'd264, 8'd231}: color_data = 12'h400;
			{9'd264, 8'd232}: color_data = 12'h900;
			{9'd264, 8'd233}: color_data = 12'ha00;
			{9'd264, 8'd234}: color_data = 12'h400;
			{9'd264, 8'd235}: color_data = 12'h310;
			{9'd264, 8'd236}: color_data = 12'hc30;
			{9'd264, 8'd237}: color_data = 12'hc20;
			{9'd264, 8'd238}: color_data = 12'h600;
			{9'd264, 8'd239}: color_data = 12'h000;
			{9'd265, 8'd68}: color_data = 12'h047;
			{9'd265, 8'd69}: color_data = 12'h6df;
			{9'd265, 8'd70}: color_data = 12'hfff;
			{9'd265, 8'd71}: color_data = 12'hcbb;
			{9'd265, 8'd72}: color_data = 12'h323;
			{9'd265, 8'd73}: color_data = 12'h002;
			{9'd265, 8'd74}: color_data = 12'h000;
			{9'd265, 8'd75}: color_data = 12'h012;
			{9'd265, 8'd76}: color_data = 12'h08c;
			{9'd265, 8'd77}: color_data = 12'h034;
			{9'd265, 8'd170}: color_data = 12'h000;
			{9'd265, 8'd171}: color_data = 12'h068;
			{9'd265, 8'd172}: color_data = 12'h8ef;
			{9'd265, 8'd173}: color_data = 12'hfff;
			{9'd265, 8'd174}: color_data = 12'haa9;
			{9'd265, 8'd175}: color_data = 12'h213;
			{9'd265, 8'd176}: color_data = 12'h002;
			{9'd265, 8'd178}: color_data = 12'h023;
			{9'd265, 8'd179}: color_data = 12'h08c;
			{9'd265, 8'd180}: color_data = 12'h023;
			{9'd265, 8'd222}: color_data = 12'h200;
			{9'd265, 8'd223}: color_data = 12'h900;
			{9'd265, 8'd224}: color_data = 12'ha00;
			{9'd265, 8'd225}: color_data = 12'h800;
			{9'd265, 8'd226}: color_data = 12'h100;
			{9'd265, 8'd227}: color_data = 12'h100;
			{9'd265, 8'd228}: color_data = 12'h300;
			{9'd265, 8'd229}: color_data = 12'h200;
			{9'd265, 8'd230}: color_data = 12'h000;
			{9'd265, 8'd231}: color_data = 12'h500;
			{9'd265, 8'd232}: color_data = 12'ha00;
			{9'd265, 8'd233}: color_data = 12'ha00;
			{9'd265, 8'd234}: color_data = 12'h500;
			{9'd265, 8'd235}: color_data = 12'h000;
			{9'd265, 8'd236}: color_data = 12'h200;
			{9'd265, 8'd237}: color_data = 12'h300;
			{9'd265, 8'd238}: color_data = 12'h100;
			{9'd265, 8'd239}: color_data = 12'h000;
			{9'd266, 8'd68}: color_data = 12'h047;
			{9'd266, 8'd69}: color_data = 12'h6ef;
			{9'd266, 8'd70}: color_data = 12'hddc;
			{9'd266, 8'd71}: color_data = 12'h434;
			{9'd266, 8'd72}: color_data = 12'h003;
			{9'd266, 8'd73}: color_data = 12'h005;
			{9'd266, 8'd74}: color_data = 12'h002;
			{9'd266, 8'd75}: color_data = 12'h012;
			{9'd266, 8'd76}: color_data = 12'h08c;
			{9'd266, 8'd77}: color_data = 12'h034;
			{9'd266, 8'd170}: color_data = 12'h000;
			{9'd266, 8'd171}: color_data = 12'h068;
			{9'd266, 8'd172}: color_data = 12'h8ff;
			{9'd266, 8'd173}: color_data = 12'hcbb;
			{9'd266, 8'd174}: color_data = 12'h223;
			{9'd266, 8'd175}: color_data = 12'h003;
			{9'd266, 8'd176}: color_data = 12'h005;
			{9'd266, 8'd177}: color_data = 12'h002;
			{9'd266, 8'd178}: color_data = 12'h023;
			{9'd266, 8'd179}: color_data = 12'h09c;
			{9'd266, 8'd180}: color_data = 12'h023;
			{9'd266, 8'd222}: color_data = 12'h300;
			{9'd266, 8'd223}: color_data = 12'hc20;
			{9'd266, 8'd224}: color_data = 12'ha00;
			{9'd266, 8'd225}: color_data = 12'h800;
			{9'd266, 8'd226}: color_data = 12'h100;
			{9'd266, 8'd227}: color_data = 12'h300;
			{9'd266, 8'd228}: color_data = 12'h500;
			{9'd266, 8'd229}: color_data = 12'h500;
			{9'd266, 8'd230}: color_data = 12'h100;
			{9'd266, 8'd231}: color_data = 12'h710;
			{9'd266, 8'd232}: color_data = 12'hc10;
			{9'd266, 8'd233}: color_data = 12'h900;
			{9'd266, 8'd234}: color_data = 12'h500;
			{9'd266, 8'd235}: color_data = 12'h100;
			{9'd266, 8'd236}: color_data = 12'h500;
			{9'd266, 8'd237}: color_data = 12'h600;
			{9'd266, 8'd238}: color_data = 12'h400;
			{9'd266, 8'd239}: color_data = 12'h000;
			{9'd267, 8'd68}: color_data = 12'h057;
			{9'd267, 8'd69}: color_data = 12'h3bd;
			{9'd267, 8'd70}: color_data = 12'h555;
			{9'd267, 8'd71}: color_data = 12'h002;
			{9'd267, 8'd72}: color_data = 12'h005;
			{9'd267, 8'd73}: color_data = 12'h005;
			{9'd267, 8'd74}: color_data = 12'h004;
			{9'd267, 8'd75}: color_data = 12'h025;
			{9'd267, 8'd76}: color_data = 12'h09c;
			{9'd267, 8'd77}: color_data = 12'h034;
			{9'd267, 8'd170}: color_data = 12'h000;
			{9'd267, 8'd171}: color_data = 12'h079;
			{9'd267, 8'd172}: color_data = 12'h4bd;
			{9'd267, 8'd173}: color_data = 12'h444;
			{9'd267, 8'd174}: color_data = 12'h002;
			{9'd267, 8'd175}: color_data = 12'h005;
			{9'd267, 8'd176}: color_data = 12'h005;
			{9'd267, 8'd177}: color_data = 12'h004;
			{9'd267, 8'd178}: color_data = 12'h036;
			{9'd267, 8'd179}: color_data = 12'h09c;
			{9'd267, 8'd180}: color_data = 12'h023;
			{9'd267, 8'd222}: color_data = 12'h410;
			{9'd267, 8'd223}: color_data = 12'hd30;
			{9'd267, 8'd224}: color_data = 12'hb00;
			{9'd267, 8'd225}: color_data = 12'h700;
			{9'd267, 8'd226}: color_data = 12'h200;
			{9'd267, 8'd227}: color_data = 12'h700;
			{9'd267, 8'd228}: color_data = 12'hb00;
			{9'd267, 8'd229}: color_data = 12'ha00;
			{9'd267, 8'd230}: color_data = 12'h300;
			{9'd267, 8'd231}: color_data = 12'h820;
			{9'd267, 8'd232}: color_data = 12'hd20;
			{9'd267, 8'd233}: color_data = 12'h900;
			{9'd267, 8'd234}: color_data = 12'h500;
			{9'd267, 8'd235}: color_data = 12'h300;
			{9'd267, 8'd236}: color_data = 12'h900;
			{9'd267, 8'd237}: color_data = 12'hb00;
			{9'd267, 8'd238}: color_data = 12'h800;
			{9'd267, 8'd239}: color_data = 12'h100;
			{9'd268, 8'd68}: color_data = 12'h036;
			{9'd268, 8'd69}: color_data = 12'h047;
			{9'd268, 8'd70}: color_data = 12'h001;
			{9'd268, 8'd71}: color_data = 12'h004;
			{9'd268, 8'd72}: color_data = 12'h004;
			{9'd268, 8'd73}: color_data = 12'h004;
			{9'd268, 8'd74}: color_data = 12'h004;
			{9'd268, 8'd75}: color_data = 12'h015;
			{9'd268, 8'd76}: color_data = 12'h059;
			{9'd268, 8'd77}: color_data = 12'h023;
			{9'd268, 8'd170}: color_data = 12'h000;
			{9'd268, 8'd171}: color_data = 12'h047;
			{9'd268, 8'd172}: color_data = 12'h036;
			{9'd268, 8'd173}: color_data = 12'h001;
			{9'd268, 8'd174}: color_data = 12'h004;
			{9'd268, 8'd175}: color_data = 12'h004;
			{9'd268, 8'd176}: color_data = 12'h004;
			{9'd268, 8'd177}: color_data = 12'h004;
			{9'd268, 8'd178}: color_data = 12'h016;
			{9'd268, 8'd179}: color_data = 12'h059;
			{9'd268, 8'd180}: color_data = 12'h012;
			{9'd268, 8'd222}: color_data = 12'h410;
			{9'd268, 8'd223}: color_data = 12'he40;
			{9'd268, 8'd224}: color_data = 12'hd20;
			{9'd268, 8'd225}: color_data = 12'h800;
			{9'd268, 8'd226}: color_data = 12'h200;
			{9'd268, 8'd227}: color_data = 12'h600;
			{9'd268, 8'd228}: color_data = 12'ha00;
			{9'd268, 8'd229}: color_data = 12'h900;
			{9'd268, 8'd230}: color_data = 12'h300;
			{9'd268, 8'd231}: color_data = 12'h820;
			{9'd268, 8'd232}: color_data = 12'hf30;
			{9'd268, 8'd233}: color_data = 12'hc00;
			{9'd268, 8'd234}: color_data = 12'h500;
			{9'd268, 8'd235}: color_data = 12'h200;
			{9'd268, 8'd236}: color_data = 12'h900;
			{9'd268, 8'd237}: color_data = 12'ha00;
			{9'd268, 8'd238}: color_data = 12'h700;
			{9'd268, 8'd239}: color_data = 12'h100;
			{9'd269, 8'd68}: color_data = 12'h013;
			{9'd269, 8'd69}: color_data = 12'h027;
			{9'd269, 8'd70}: color_data = 12'h016;
			{9'd269, 8'd71}: color_data = 12'h027;
			{9'd269, 8'd72}: color_data = 12'h027;
			{9'd269, 8'd73}: color_data = 12'h017;
			{9'd269, 8'd74}: color_data = 12'h027;
			{9'd269, 8'd75}: color_data = 12'h028;
			{9'd269, 8'd76}: color_data = 12'h027;
			{9'd269, 8'd77}: color_data = 12'h001;
			{9'd269, 8'd170}: color_data = 12'h000;
			{9'd269, 8'd171}: color_data = 12'h014;
			{9'd269, 8'd172}: color_data = 12'h027;
			{9'd269, 8'd173}: color_data = 12'h016;
			{9'd269, 8'd174}: color_data = 12'h027;
			{9'd269, 8'd175}: color_data = 12'h027;
			{9'd269, 8'd176}: color_data = 12'h017;
			{9'd269, 8'd177}: color_data = 12'h027;
			{9'd269, 8'd178}: color_data = 12'h028;
			{9'd269, 8'd179}: color_data = 12'h026;
			{9'd269, 8'd180}: color_data = 12'h001;
			{9'd269, 8'd222}: color_data = 12'h300;
			{9'd269, 8'd223}: color_data = 12'hc30;
			{9'd269, 8'd224}: color_data = 12'hc30;
			{9'd269, 8'd225}: color_data = 12'h600;
			{9'd269, 8'd226}: color_data = 12'h100;
			{9'd269, 8'd227}: color_data = 12'h600;
			{9'd269, 8'd228}: color_data = 12'ha00;
			{9'd269, 8'd229}: color_data = 12'h900;
			{9'd269, 8'd230}: color_data = 12'h300;
			{9'd269, 8'd231}: color_data = 12'h620;
			{9'd269, 8'd232}: color_data = 12'hd40;
			{9'd269, 8'd233}: color_data = 12'ha20;
			{9'd269, 8'd234}: color_data = 12'h300;
			{9'd269, 8'd235}: color_data = 12'h200;
			{9'd269, 8'd236}: color_data = 12'h900;
			{9'd269, 8'd237}: color_data = 12'ha00;
			{9'd269, 8'd238}: color_data = 12'h700;
			{9'd269, 8'd239}: color_data = 12'h100;
			{9'd270, 8'd68}: color_data = 12'h045;
			{9'd270, 8'd69}: color_data = 12'h09e;
			{9'd270, 8'd70}: color_data = 12'h09e;
			{9'd270, 8'd71}: color_data = 12'h09e;
			{9'd270, 8'd72}: color_data = 12'h09e;
			{9'd270, 8'd73}: color_data = 12'h09e;
			{9'd270, 8'd74}: color_data = 12'h09e;
			{9'd270, 8'd75}: color_data = 12'h09e;
			{9'd270, 8'd76}: color_data = 12'h08c;
			{9'd270, 8'd77}: color_data = 12'h023;
			{9'd270, 8'd170}: color_data = 12'h000;
			{9'd270, 8'd171}: color_data = 12'h057;
			{9'd270, 8'd172}: color_data = 12'h0ae;
			{9'd270, 8'd173}: color_data = 12'h09e;
			{9'd270, 8'd174}: color_data = 12'h09e;
			{9'd270, 8'd175}: color_data = 12'h09e;
			{9'd270, 8'd176}: color_data = 12'h09e;
			{9'd270, 8'd177}: color_data = 12'h09e;
			{9'd270, 8'd178}: color_data = 12'h09e;
			{9'd270, 8'd179}: color_data = 12'h07b;
			{9'd270, 8'd180}: color_data = 12'h012;
			{9'd270, 8'd222}: color_data = 12'h000;
			{9'd270, 8'd223}: color_data = 12'h200;
			{9'd270, 8'd224}: color_data = 12'h300;
			{9'd270, 8'd225}: color_data = 12'h100;
			{9'd270, 8'd226}: color_data = 12'h000;
			{9'd270, 8'd227}: color_data = 12'h700;
			{9'd270, 8'd228}: color_data = 12'ha00;
			{9'd270, 8'd229}: color_data = 12'h900;
			{9'd270, 8'd230}: color_data = 12'h300;
			{9'd270, 8'd231}: color_data = 12'h000;
			{9'd270, 8'd232}: color_data = 12'h310;
			{9'd270, 8'd233}: color_data = 12'h200;
			{9'd270, 8'd234}: color_data = 12'h000;
			{9'd270, 8'd235}: color_data = 12'h300;
			{9'd270, 8'd236}: color_data = 12'h900;
			{9'd270, 8'd237}: color_data = 12'ha00;
			{9'd270, 8'd238}: color_data = 12'h700;
			{9'd270, 8'd239}: color_data = 12'h100;
			{9'd271, 8'd68}: color_data = 12'h057;
			{9'd271, 8'd69}: color_data = 12'h4ef;
			{9'd271, 8'd70}: color_data = 12'h7ef;
			{9'd271, 8'd71}: color_data = 12'h0cf;
			{9'd271, 8'd72}: color_data = 12'h0cf;
			{9'd271, 8'd73}: color_data = 12'h0df;
			{9'd271, 8'd74}: color_data = 12'h0bd;
			{9'd271, 8'd75}: color_data = 12'h068;
			{9'd271, 8'd76}: color_data = 12'h09c;
			{9'd271, 8'd77}: color_data = 12'h034;
			{9'd271, 8'd170}: color_data = 12'h000;
			{9'd271, 8'd171}: color_data = 12'h069;
			{9'd271, 8'd172}: color_data = 12'h6ef;
			{9'd271, 8'd173}: color_data = 12'h6ef;
			{9'd271, 8'd174}: color_data = 12'h0cf;
			{9'd271, 8'd175}: color_data = 12'h0cf;
			{9'd271, 8'd176}: color_data = 12'h0df;
			{9'd271, 8'd177}: color_data = 12'h0ac;
			{9'd271, 8'd178}: color_data = 12'h079;
			{9'd271, 8'd179}: color_data = 12'h09c;
			{9'd271, 8'd180}: color_data = 12'h023;
			{9'd271, 8'd222}: color_data = 12'h100;
			{9'd271, 8'd223}: color_data = 12'h400;
			{9'd271, 8'd224}: color_data = 12'h500;
			{9'd271, 8'd225}: color_data = 12'h400;
			{9'd271, 8'd226}: color_data = 12'h200;
			{9'd271, 8'd227}: color_data = 12'ha20;
			{9'd271, 8'd228}: color_data = 12'hb10;
			{9'd271, 8'd229}: color_data = 12'h900;
			{9'd271, 8'd230}: color_data = 12'h300;
			{9'd271, 8'd231}: color_data = 12'h200;
			{9'd271, 8'd232}: color_data = 12'h500;
			{9'd271, 8'd233}: color_data = 12'h500;
			{9'd271, 8'd234}: color_data = 12'h200;
			{9'd271, 8'd235}: color_data = 12'h410;
			{9'd271, 8'd236}: color_data = 12'hc20;
			{9'd271, 8'd237}: color_data = 12'ha00;
			{9'd271, 8'd238}: color_data = 12'h700;
			{9'd271, 8'd239}: color_data = 12'h100;
			{9'd272, 8'd68}: color_data = 12'h047;
			{9'd272, 8'd69}: color_data = 12'h6df;
			{9'd272, 8'd70}: color_data = 12'heff;
			{9'd272, 8'd71}: color_data = 12'h6df;
			{9'd272, 8'd72}: color_data = 12'h0bf;
			{9'd272, 8'd73}: color_data = 12'h0be;
			{9'd272, 8'd74}: color_data = 12'h056;
			{9'd272, 8'd75}: color_data = 12'h012;
			{9'd272, 8'd76}: color_data = 12'h08b;
			{9'd272, 8'd77}: color_data = 12'h034;
			{9'd272, 8'd170}: color_data = 12'h000;
			{9'd272, 8'd171}: color_data = 12'h068;
			{9'd272, 8'd172}: color_data = 12'h8ef;
			{9'd272, 8'd173}: color_data = 12'hdff;
			{9'd272, 8'd174}: color_data = 12'h4cf;
			{9'd272, 8'd175}: color_data = 12'h0cf;
			{9'd272, 8'd176}: color_data = 12'h0ae;
			{9'd272, 8'd177}: color_data = 12'h035;
			{9'd272, 8'd178}: color_data = 12'h023;
			{9'd272, 8'd179}: color_data = 12'h08c;
			{9'd272, 8'd180}: color_data = 12'h023;
			{9'd272, 8'd222}: color_data = 12'h200;
			{9'd272, 8'd223}: color_data = 12'h900;
			{9'd272, 8'd224}: color_data = 12'hb00;
			{9'd272, 8'd225}: color_data = 12'h800;
			{9'd272, 8'd226}: color_data = 12'h200;
			{9'd272, 8'd227}: color_data = 12'hb30;
			{9'd272, 8'd228}: color_data = 12'hc10;
			{9'd272, 8'd229}: color_data = 12'h800;
			{9'd272, 8'd230}: color_data = 12'h300;
			{9'd272, 8'd231}: color_data = 12'h500;
			{9'd272, 8'd232}: color_data = 12'ha00;
			{9'd272, 8'd233}: color_data = 12'ha00;
			{9'd272, 8'd234}: color_data = 12'h500;
			{9'd272, 8'd235}: color_data = 12'h510;
			{9'd272, 8'd236}: color_data = 12'hd30;
			{9'd272, 8'd237}: color_data = 12'ha00;
			{9'd272, 8'd238}: color_data = 12'h700;
			{9'd272, 8'd239}: color_data = 12'h100;
			{9'd273, 8'd68}: color_data = 12'h047;
			{9'd273, 8'd69}: color_data = 12'h6df;
			{9'd273, 8'd70}: color_data = 12'hfff;
			{9'd273, 8'd71}: color_data = 12'hdff;
			{9'd273, 8'd72}: color_data = 12'h5df;
			{9'd273, 8'd73}: color_data = 12'h068;
			{9'd273, 8'd74}: color_data = 12'h000;
			{9'd273, 8'd75}: color_data = 12'h012;
			{9'd273, 8'd76}: color_data = 12'h08c;
			{9'd273, 8'd77}: color_data = 12'h034;
			{9'd273, 8'd170}: color_data = 12'h000;
			{9'd273, 8'd171}: color_data = 12'h068;
			{9'd273, 8'd172}: color_data = 12'h8ef;
			{9'd273, 8'd173}: color_data = 12'hfff;
			{9'd273, 8'd174}: color_data = 12'hcff;
			{9'd273, 8'd175}: color_data = 12'h4ce;
			{9'd273, 8'd176}: color_data = 12'h057;
			{9'd273, 8'd177}: color_data = 12'h000;
			{9'd273, 8'd178}: color_data = 12'h023;
			{9'd273, 8'd179}: color_data = 12'h08c;
			{9'd273, 8'd180}: color_data = 12'h023;
			{9'd273, 8'd222}: color_data = 12'h200;
			{9'd273, 8'd223}: color_data = 12'h900;
			{9'd273, 8'd224}: color_data = 12'ha00;
			{9'd273, 8'd225}: color_data = 12'h700;
			{9'd273, 8'd226}: color_data = 12'h200;
			{9'd273, 8'd227}: color_data = 12'hb30;
			{9'd273, 8'd228}: color_data = 12'he20;
			{9'd273, 8'd229}: color_data = 12'ha00;
			{9'd273, 8'd230}: color_data = 12'h300;
			{9'd273, 8'd231}: color_data = 12'h400;
			{9'd273, 8'd232}: color_data = 12'ha00;
			{9'd273, 8'd233}: color_data = 12'ha00;
			{9'd273, 8'd234}: color_data = 12'h400;
			{9'd273, 8'd235}: color_data = 12'h510;
			{9'd273, 8'd236}: color_data = 12'hf40;
			{9'd273, 8'd237}: color_data = 12'hd10;
			{9'd273, 8'd238}: color_data = 12'h800;
			{9'd273, 8'd239}: color_data = 12'h100;
			{9'd274, 8'd68}: color_data = 12'h047;
			{9'd274, 8'd69}: color_data = 12'h6df;
			{9'd274, 8'd70}: color_data = 12'hfff;
			{9'd274, 8'd71}: color_data = 12'hfff;
			{9'd274, 8'd72}: color_data = 12'h9aa;
			{9'd274, 8'd73}: color_data = 12'h011;
			{9'd274, 8'd75}: color_data = 12'h012;
			{9'd274, 8'd76}: color_data = 12'h08c;
			{9'd274, 8'd77}: color_data = 12'h034;
			{9'd274, 8'd170}: color_data = 12'h000;
			{9'd274, 8'd171}: color_data = 12'h068;
			{9'd274, 8'd172}: color_data = 12'h7ef;
			{9'd274, 8'd173}: color_data = 12'hfff;
			{9'd274, 8'd174}: color_data = 12'hfff;
			{9'd274, 8'd175}: color_data = 12'h899;
			{9'd274, 8'd176}: color_data = 12'h001;
			{9'd274, 8'd178}: color_data = 12'h024;
			{9'd274, 8'd179}: color_data = 12'h08c;
			{9'd274, 8'd180}: color_data = 12'h023;
			{9'd274, 8'd222}: color_data = 12'h200;
			{9'd274, 8'd223}: color_data = 12'h800;
			{9'd274, 8'd224}: color_data = 12'ha00;
			{9'd274, 8'd225}: color_data = 12'h800;
			{9'd274, 8'd226}: color_data = 12'h200;
			{9'd274, 8'd227}: color_data = 12'h920;
			{9'd274, 8'd228}: color_data = 12'hd30;
			{9'd274, 8'd229}: color_data = 12'h910;
			{9'd274, 8'd230}: color_data = 12'h200;
			{9'd274, 8'd231}: color_data = 12'h400;
			{9'd274, 8'd232}: color_data = 12'h900;
			{9'd274, 8'd233}: color_data = 12'ha00;
			{9'd274, 8'd234}: color_data = 12'h400;
			{9'd274, 8'd235}: color_data = 12'h310;
			{9'd274, 8'd236}: color_data = 12'hc30;
			{9'd274, 8'd237}: color_data = 12'hc20;
			{9'd274, 8'd238}: color_data = 12'h600;
			{9'd274, 8'd239}: color_data = 12'h000;
			{9'd275, 8'd68}: color_data = 12'h047;
			{9'd275, 8'd69}: color_data = 12'h6df;
			{9'd275, 8'd70}: color_data = 12'hfff;
			{9'd275, 8'd71}: color_data = 12'hcbb;
			{9'd275, 8'd72}: color_data = 12'h323;
			{9'd275, 8'd73}: color_data = 12'h002;
			{9'd275, 8'd74}: color_data = 12'h000;
			{9'd275, 8'd75}: color_data = 12'h012;
			{9'd275, 8'd76}: color_data = 12'h08c;
			{9'd275, 8'd77}: color_data = 12'h034;
			{9'd275, 8'd170}: color_data = 12'h000;
			{9'd275, 8'd171}: color_data = 12'h068;
			{9'd275, 8'd172}: color_data = 12'h8ef;
			{9'd275, 8'd173}: color_data = 12'hfff;
			{9'd275, 8'd174}: color_data = 12'haa9;
			{9'd275, 8'd175}: color_data = 12'h212;
			{9'd275, 8'd176}: color_data = 12'h002;
			{9'd275, 8'd177}: color_data = 12'h000;
			{9'd275, 8'd178}: color_data = 12'h023;
			{9'd275, 8'd179}: color_data = 12'h08c;
			{9'd275, 8'd180}: color_data = 12'h023;
			{9'd275, 8'd222}: color_data = 12'h200;
			{9'd275, 8'd223}: color_data = 12'h900;
			{9'd275, 8'd224}: color_data = 12'ha00;
			{9'd275, 8'd225}: color_data = 12'h800;
			{9'd275, 8'd226}: color_data = 12'h100;
			{9'd275, 8'd227}: color_data = 12'h100;
			{9'd275, 8'd228}: color_data = 12'h310;
			{9'd275, 8'd229}: color_data = 12'h200;
			{9'd275, 8'd230}: color_data = 12'h000;
			{9'd275, 8'd231}: color_data = 12'h500;
			{9'd275, 8'd232}: color_data = 12'ha00;
			{9'd275, 8'd233}: color_data = 12'ha00;
			{9'd275, 8'd234}: color_data = 12'h500;
			{9'd275, 8'd235}: color_data = 12'h000;
			{9'd275, 8'd236}: color_data = 12'h200;
			{9'd275, 8'd237}: color_data = 12'h300;
			{9'd275, 8'd238}: color_data = 12'h100;
			{9'd275, 8'd239}: color_data = 12'h000;
			{9'd276, 8'd68}: color_data = 12'h047;
			{9'd276, 8'd69}: color_data = 12'h6ef;
			{9'd276, 8'd70}: color_data = 12'hdcc;
			{9'd276, 8'd71}: color_data = 12'h433;
			{9'd276, 8'd72}: color_data = 12'h003;
			{9'd276, 8'd73}: color_data = 12'h005;
			{9'd276, 8'd74}: color_data = 12'h002;
			{9'd276, 8'd75}: color_data = 12'h012;
			{9'd276, 8'd76}: color_data = 12'h08c;
			{9'd276, 8'd77}: color_data = 12'h034;
			{9'd276, 8'd170}: color_data = 12'h000;
			{9'd276, 8'd171}: color_data = 12'h068;
			{9'd276, 8'd172}: color_data = 12'h8ff;
			{9'd276, 8'd173}: color_data = 12'hcbb;
			{9'd276, 8'd174}: color_data = 12'h323;
			{9'd276, 8'd175}: color_data = 12'h003;
			{9'd276, 8'd176}: color_data = 12'h005;
			{9'd276, 8'd177}: color_data = 12'h002;
			{9'd276, 8'd178}: color_data = 12'h023;
			{9'd276, 8'd179}: color_data = 12'h09c;
			{9'd276, 8'd180}: color_data = 12'h023;
			{9'd276, 8'd222}: color_data = 12'h300;
			{9'd276, 8'd223}: color_data = 12'hc20;
			{9'd276, 8'd224}: color_data = 12'ha00;
			{9'd276, 8'd225}: color_data = 12'h800;
			{9'd276, 8'd226}: color_data = 12'h100;
			{9'd276, 8'd227}: color_data = 12'h300;
			{9'd276, 8'd228}: color_data = 12'h500;
			{9'd276, 8'd229}: color_data = 12'h500;
			{9'd276, 8'd230}: color_data = 12'h100;
			{9'd276, 8'd231}: color_data = 12'h710;
			{9'd276, 8'd232}: color_data = 12'hc10;
			{9'd276, 8'd233}: color_data = 12'h900;
			{9'd276, 8'd234}: color_data = 12'h500;
			{9'd276, 8'd235}: color_data = 12'h100;
			{9'd276, 8'd236}: color_data = 12'h500;
			{9'd276, 8'd237}: color_data = 12'h600;
			{9'd276, 8'd238}: color_data = 12'h400;
			{9'd276, 8'd239}: color_data = 12'h000;
			{9'd277, 8'd68}: color_data = 12'h057;
			{9'd277, 8'd69}: color_data = 12'h3bd;
			{9'd277, 8'd70}: color_data = 12'h555;
			{9'd277, 8'd71}: color_data = 12'h002;
			{9'd277, 8'd72}: color_data = 12'h005;
			{9'd277, 8'd73}: color_data = 12'h005;
			{9'd277, 8'd74}: color_data = 12'h004;
			{9'd277, 8'd75}: color_data = 12'h025;
			{9'd277, 8'd76}: color_data = 12'h09c;
			{9'd277, 8'd77}: color_data = 12'h034;
			{9'd277, 8'd170}: color_data = 12'h000;
			{9'd277, 8'd171}: color_data = 12'h079;
			{9'd277, 8'd172}: color_data = 12'h4bd;
			{9'd277, 8'd173}: color_data = 12'h444;
			{9'd277, 8'd174}: color_data = 12'h002;
			{9'd277, 8'd175}: color_data = 12'h005;
			{9'd277, 8'd176}: color_data = 12'h005;
			{9'd277, 8'd177}: color_data = 12'h004;
			{9'd277, 8'd178}: color_data = 12'h036;
			{9'd277, 8'd179}: color_data = 12'h09c;
			{9'd277, 8'd180}: color_data = 12'h023;
			{9'd277, 8'd222}: color_data = 12'h410;
			{9'd277, 8'd223}: color_data = 12'hd30;
			{9'd277, 8'd224}: color_data = 12'hb00;
			{9'd277, 8'd225}: color_data = 12'h700;
			{9'd277, 8'd226}: color_data = 12'h200;
			{9'd277, 8'd227}: color_data = 12'h700;
			{9'd277, 8'd228}: color_data = 12'hb00;
			{9'd277, 8'd229}: color_data = 12'ha00;
			{9'd277, 8'd230}: color_data = 12'h300;
			{9'd277, 8'd231}: color_data = 12'h820;
			{9'd277, 8'd232}: color_data = 12'hd20;
			{9'd277, 8'd233}: color_data = 12'h900;
			{9'd277, 8'd234}: color_data = 12'h500;
			{9'd277, 8'd235}: color_data = 12'h300;
			{9'd277, 8'd236}: color_data = 12'h900;
			{9'd277, 8'd237}: color_data = 12'hb00;
			{9'd277, 8'd238}: color_data = 12'h800;
			{9'd277, 8'd239}: color_data = 12'h100;
			{9'd278, 8'd68}: color_data = 12'h035;
			{9'd278, 8'd69}: color_data = 12'h047;
			{9'd278, 8'd70}: color_data = 12'h001;
			{9'd278, 8'd71}: color_data = 12'h004;
			{9'd278, 8'd72}: color_data = 12'h004;
			{9'd278, 8'd73}: color_data = 12'h004;
			{9'd278, 8'd74}: color_data = 12'h004;
			{9'd278, 8'd75}: color_data = 12'h015;
			{9'd278, 8'd76}: color_data = 12'h059;
			{9'd278, 8'd77}: color_data = 12'h023;
			{9'd278, 8'd170}: color_data = 12'h000;
			{9'd278, 8'd171}: color_data = 12'h047;
			{9'd278, 8'd172}: color_data = 12'h036;
			{9'd278, 8'd173}: color_data = 12'h001;
			{9'd278, 8'd174}: color_data = 12'h004;
			{9'd278, 8'd175}: color_data = 12'h004;
			{9'd278, 8'd176}: color_data = 12'h004;
			{9'd278, 8'd177}: color_data = 12'h004;
			{9'd278, 8'd178}: color_data = 12'h016;
			{9'd278, 8'd179}: color_data = 12'h059;
			{9'd278, 8'd180}: color_data = 12'h012;
			{9'd278, 8'd222}: color_data = 12'h410;
			{9'd278, 8'd223}: color_data = 12'he40;
			{9'd278, 8'd224}: color_data = 12'hd20;
			{9'd278, 8'd225}: color_data = 12'h800;
			{9'd278, 8'd226}: color_data = 12'h200;
			{9'd278, 8'd227}: color_data = 12'h600;
			{9'd278, 8'd228}: color_data = 12'ha00;
			{9'd278, 8'd229}: color_data = 12'h900;
			{9'd278, 8'd230}: color_data = 12'h300;
			{9'd278, 8'd231}: color_data = 12'h820;
			{9'd278, 8'd232}: color_data = 12'hf30;
			{9'd278, 8'd233}: color_data = 12'hc00;
			{9'd278, 8'd234}: color_data = 12'h500;
			{9'd278, 8'd235}: color_data = 12'h200;
			{9'd278, 8'd236}: color_data = 12'h900;
			{9'd278, 8'd237}: color_data = 12'ha00;
			{9'd278, 8'd238}: color_data = 12'h700;
			{9'd278, 8'd239}: color_data = 12'h100;
			{9'd279, 8'd15}: color_data = 12'h000;
			{9'd279, 8'd16}: color_data = 12'h110;
			{9'd279, 8'd17}: color_data = 12'h332;
			{9'd279, 8'd18}: color_data = 12'h333;
			{9'd279, 8'd19}: color_data = 12'h222;
			{9'd279, 8'd20}: color_data = 12'h333;
			{9'd279, 8'd21}: color_data = 12'h221;
			{9'd279, 8'd22}: color_data = 12'h120;
			{9'd279, 8'd23}: color_data = 12'h120;
			{9'd279, 8'd24}: color_data = 12'h120;
			{9'd279, 8'd25}: color_data = 12'h120;
			{9'd279, 8'd26}: color_data = 12'h110;
			{9'd279, 8'd27}: color_data = 12'h010;
			{9'd279, 8'd28}: color_data = 12'h000;
			{9'd279, 8'd29}: color_data = 12'h000;
			{9'd279, 8'd30}: color_data = 12'h000;
			{9'd279, 8'd31}: color_data = 12'h110;
			{9'd279, 8'd32}: color_data = 12'h110;
			{9'd279, 8'd33}: color_data = 12'h000;
			{9'd279, 8'd68}: color_data = 12'h013;
			{9'd279, 8'd69}: color_data = 12'h027;
			{9'd279, 8'd70}: color_data = 12'h016;
			{9'd279, 8'd71}: color_data = 12'h027;
			{9'd279, 8'd72}: color_data = 12'h027;
			{9'd279, 8'd73}: color_data = 12'h027;
			{9'd279, 8'd74}: color_data = 12'h027;
			{9'd279, 8'd75}: color_data = 12'h028;
			{9'd279, 8'd76}: color_data = 12'h027;
			{9'd279, 8'd77}: color_data = 12'h001;
			{9'd279, 8'd128}: color_data = 12'h001;
			{9'd279, 8'd129}: color_data = 12'h023;
			{9'd279, 8'd130}: color_data = 12'h012;
			{9'd279, 8'd131}: color_data = 12'h022;
			{9'd279, 8'd132}: color_data = 12'h022;
			{9'd279, 8'd133}: color_data = 12'h022;
			{9'd279, 8'd134}: color_data = 12'h023;
			{9'd279, 8'd135}: color_data = 12'h023;
			{9'd279, 8'd136}: color_data = 12'h022;
			{9'd279, 8'd137}: color_data = 12'h000;
			{9'd279, 8'd170}: color_data = 12'h000;
			{9'd279, 8'd171}: color_data = 12'h014;
			{9'd279, 8'd172}: color_data = 12'h027;
			{9'd279, 8'd173}: color_data = 12'h016;
			{9'd279, 8'd174}: color_data = 12'h027;
			{9'd279, 8'd175}: color_data = 12'h027;
			{9'd279, 8'd176}: color_data = 12'h027;
			{9'd279, 8'd177}: color_data = 12'h027;
			{9'd279, 8'd178}: color_data = 12'h028;
			{9'd279, 8'd179}: color_data = 12'h026;
			{9'd279, 8'd180}: color_data = 12'h001;
			{9'd279, 8'd222}: color_data = 12'h300;
			{9'd279, 8'd223}: color_data = 12'hc30;
			{9'd279, 8'd224}: color_data = 12'hc30;
			{9'd279, 8'd225}: color_data = 12'h600;
			{9'd279, 8'd226}: color_data = 12'h100;
			{9'd279, 8'd227}: color_data = 12'h600;
			{9'd279, 8'd228}: color_data = 12'ha00;
			{9'd279, 8'd229}: color_data = 12'h900;
			{9'd279, 8'd230}: color_data = 12'h300;
			{9'd279, 8'd231}: color_data = 12'h620;
			{9'd279, 8'd232}: color_data = 12'hd40;
			{9'd279, 8'd233}: color_data = 12'ha20;
			{9'd279, 8'd234}: color_data = 12'h300;
			{9'd279, 8'd235}: color_data = 12'h200;
			{9'd279, 8'd236}: color_data = 12'h900;
			{9'd279, 8'd237}: color_data = 12'ha00;
			{9'd279, 8'd238}: color_data = 12'h700;
			{9'd279, 8'd239}: color_data = 12'h100;
			{9'd280, 8'd15}: color_data = 12'h010;
			{9'd280, 8'd16}: color_data = 12'h681;
			{9'd280, 8'd17}: color_data = 12'hcd9;
			{9'd280, 8'd18}: color_data = 12'hddd;
			{9'd280, 8'd19}: color_data = 12'hddd;
			{9'd280, 8'd20}: color_data = 12'hddd;
			{9'd280, 8'd21}: color_data = 12'hab5;
			{9'd280, 8'd22}: color_data = 12'h790;
			{9'd280, 8'd23}: color_data = 12'h790;
			{9'd280, 8'd24}: color_data = 12'h790;
			{9'd280, 8'd25}: color_data = 12'h890;
			{9'd280, 8'd26}: color_data = 12'h780;
			{9'd280, 8'd27}: color_data = 12'h440;
			{9'd280, 8'd28}: color_data = 12'h020;
			{9'd280, 8'd29}: color_data = 12'h130;
			{9'd280, 8'd30}: color_data = 12'h240;
			{9'd280, 8'd31}: color_data = 12'h550;
			{9'd280, 8'd32}: color_data = 12'h550;
			{9'd280, 8'd33}: color_data = 12'h110;
			{9'd280, 8'd68}: color_data = 12'h035;
			{9'd280, 8'd69}: color_data = 12'h09e;
			{9'd280, 8'd70}: color_data = 12'h09e;
			{9'd280, 8'd71}: color_data = 12'h09e;
			{9'd280, 8'd72}: color_data = 12'h09e;
			{9'd280, 8'd73}: color_data = 12'h09e;
			{9'd280, 8'd74}: color_data = 12'h09e;
			{9'd280, 8'd75}: color_data = 12'h09e;
			{9'd280, 8'd76}: color_data = 12'h08c;
			{9'd280, 8'd77}: color_data = 12'h023;
			{9'd280, 8'd128}: color_data = 12'h045;
			{9'd280, 8'd129}: color_data = 12'h0ad;
			{9'd280, 8'd130}: color_data = 12'h09d;
			{9'd280, 8'd131}: color_data = 12'h09d;
			{9'd280, 8'd132}: color_data = 12'h09d;
			{9'd280, 8'd133}: color_data = 12'h09d;
			{9'd280, 8'd134}: color_data = 12'h09d;
			{9'd280, 8'd135}: color_data = 12'h09d;
			{9'd280, 8'd136}: color_data = 12'h09c;
			{9'd280, 8'd137}: color_data = 12'h023;
			{9'd280, 8'd170}: color_data = 12'h000;
			{9'd280, 8'd171}: color_data = 12'h057;
			{9'd280, 8'd172}: color_data = 12'h0ae;
			{9'd280, 8'd173}: color_data = 12'h09e;
			{9'd280, 8'd174}: color_data = 12'h09e;
			{9'd280, 8'd175}: color_data = 12'h09e;
			{9'd280, 8'd176}: color_data = 12'h09e;
			{9'd280, 8'd177}: color_data = 12'h09e;
			{9'd280, 8'd178}: color_data = 12'h09e;
			{9'd280, 8'd179}: color_data = 12'h07b;
			{9'd280, 8'd180}: color_data = 12'h012;
			{9'd280, 8'd222}: color_data = 12'h000;
			{9'd280, 8'd223}: color_data = 12'h200;
			{9'd280, 8'd224}: color_data = 12'h300;
			{9'd280, 8'd225}: color_data = 12'h100;
			{9'd280, 8'd226}: color_data = 12'h000;
			{9'd280, 8'd227}: color_data = 12'h700;
			{9'd280, 8'd228}: color_data = 12'ha00;
			{9'd280, 8'd229}: color_data = 12'h900;
			{9'd280, 8'd230}: color_data = 12'h300;
			{9'd280, 8'd231}: color_data = 12'h100;
			{9'd280, 8'd232}: color_data = 12'h310;
			{9'd280, 8'd233}: color_data = 12'h200;
			{9'd280, 8'd234}: color_data = 12'h000;
			{9'd280, 8'd235}: color_data = 12'h300;
			{9'd280, 8'd236}: color_data = 12'h900;
			{9'd280, 8'd237}: color_data = 12'ha00;
			{9'd280, 8'd238}: color_data = 12'h700;
			{9'd280, 8'd239}: color_data = 12'h100;
			{9'd281, 8'd15}: color_data = 12'h110;
			{9'd281, 8'd16}: color_data = 12'h8a0;
			{9'd281, 8'd17}: color_data = 12'hce5;
			{9'd281, 8'd18}: color_data = 12'hffd;
			{9'd281, 8'd19}: color_data = 12'hfff;
			{9'd281, 8'd20}: color_data = 12'heea;
			{9'd281, 8'd21}: color_data = 12'hbc2;
			{9'd281, 8'd22}: color_data = 12'h9c0;
			{9'd281, 8'd23}: color_data = 12'hac0;
			{9'd281, 8'd24}: color_data = 12'hac0;
			{9'd281, 8'd25}: color_data = 12'hac0;
			{9'd281, 8'd26}: color_data = 12'h9b0;
			{9'd281, 8'd27}: color_data = 12'h550;
			{9'd281, 8'd28}: color_data = 12'h020;
			{9'd281, 8'd29}: color_data = 12'h140;
			{9'd281, 8'd30}: color_data = 12'h250;
			{9'd281, 8'd31}: color_data = 12'h660;
			{9'd281, 8'd32}: color_data = 12'h760;
			{9'd281, 8'd33}: color_data = 12'h110;
			{9'd281, 8'd68}: color_data = 12'h057;
			{9'd281, 8'd69}: color_data = 12'h4ef;
			{9'd281, 8'd70}: color_data = 12'h7ef;
			{9'd281, 8'd71}: color_data = 12'h0cf;
			{9'd281, 8'd72}: color_data = 12'h0cf;
			{9'd281, 8'd73}: color_data = 12'h0df;
			{9'd281, 8'd74}: color_data = 12'h0bd;
			{9'd281, 8'd75}: color_data = 12'h068;
			{9'd281, 8'd76}: color_data = 12'h09c;
			{9'd281, 8'd77}: color_data = 12'h034;
			{9'd281, 8'd128}: color_data = 12'h057;
			{9'd281, 8'd129}: color_data = 12'h4ef;
			{9'd281, 8'd130}: color_data = 12'h7ef;
			{9'd281, 8'd131}: color_data = 12'h0cf;
			{9'd281, 8'd132}: color_data = 12'h0cf;
			{9'd281, 8'd133}: color_data = 12'h0df;
			{9'd281, 8'd134}: color_data = 12'h0be;
			{9'd281, 8'd135}: color_data = 12'h069;
			{9'd281, 8'd136}: color_data = 12'h09c;
			{9'd281, 8'd137}: color_data = 12'h034;
			{9'd281, 8'd170}: color_data = 12'h000;
			{9'd281, 8'd171}: color_data = 12'h069;
			{9'd281, 8'd172}: color_data = 12'h6ef;
			{9'd281, 8'd173}: color_data = 12'h6ef;
			{9'd281, 8'd174}: color_data = 12'h0cf;
			{9'd281, 8'd175}: color_data = 12'h0cf;
			{9'd281, 8'd176}: color_data = 12'h0df;
			{9'd281, 8'd177}: color_data = 12'h0ac;
			{9'd281, 8'd178}: color_data = 12'h079;
			{9'd281, 8'd179}: color_data = 12'h09c;
			{9'd281, 8'd180}: color_data = 12'h023;
			{9'd281, 8'd222}: color_data = 12'h100;
			{9'd281, 8'd223}: color_data = 12'h500;
			{9'd281, 8'd224}: color_data = 12'h600;
			{9'd281, 8'd225}: color_data = 12'h400;
			{9'd281, 8'd226}: color_data = 12'h200;
			{9'd281, 8'd227}: color_data = 12'ha20;
			{9'd281, 8'd228}: color_data = 12'hb10;
			{9'd281, 8'd229}: color_data = 12'h900;
			{9'd281, 8'd230}: color_data = 12'h300;
			{9'd281, 8'd231}: color_data = 12'h200;
			{9'd281, 8'd232}: color_data = 12'h500;
			{9'd281, 8'd233}: color_data = 12'h500;
			{9'd281, 8'd234}: color_data = 12'h200;
			{9'd281, 8'd235}: color_data = 12'h410;
			{9'd281, 8'd236}: color_data = 12'hc20;
			{9'd281, 8'd237}: color_data = 12'ha00;
			{9'd281, 8'd238}: color_data = 12'h700;
			{9'd281, 8'd239}: color_data = 12'h100;
			{9'd282, 8'd15}: color_data = 12'h110;
			{9'd282, 8'd16}: color_data = 12'h790;
			{9'd282, 8'd17}: color_data = 12'h9c0;
			{9'd282, 8'd18}: color_data = 12'heeb;
			{9'd282, 8'd19}: color_data = 12'hfff;
			{9'd282, 8'd20}: color_data = 12'hbd6;
			{9'd282, 8'd21}: color_data = 12'h8b0;
			{9'd282, 8'd22}: color_data = 12'h9b0;
			{9'd282, 8'd23}: color_data = 12'h9b0;
			{9'd282, 8'd24}: color_data = 12'h9b0;
			{9'd282, 8'd25}: color_data = 12'h9b0;
			{9'd282, 8'd26}: color_data = 12'h9a0;
			{9'd282, 8'd27}: color_data = 12'h550;
			{9'd282, 8'd28}: color_data = 12'h020;
			{9'd282, 8'd29}: color_data = 12'h130;
			{9'd282, 8'd30}: color_data = 12'h240;
			{9'd282, 8'd31}: color_data = 12'h660;
			{9'd282, 8'd32}: color_data = 12'h660;
			{9'd282, 8'd33}: color_data = 12'h110;
			{9'd282, 8'd68}: color_data = 12'h047;
			{9'd282, 8'd69}: color_data = 12'h6df;
			{9'd282, 8'd70}: color_data = 12'heff;
			{9'd282, 8'd71}: color_data = 12'h6df;
			{9'd282, 8'd72}: color_data = 12'h0bf;
			{9'd282, 8'd73}: color_data = 12'h0be;
			{9'd282, 8'd74}: color_data = 12'h056;
			{9'd282, 8'd75}: color_data = 12'h012;
			{9'd282, 8'd76}: color_data = 12'h08b;
			{9'd282, 8'd77}: color_data = 12'h034;
			{9'd282, 8'd128}: color_data = 12'h047;
			{9'd282, 8'd129}: color_data = 12'h6df;
			{9'd282, 8'd130}: color_data = 12'heff;
			{9'd282, 8'd131}: color_data = 12'h6df;
			{9'd282, 8'd132}: color_data = 12'h0bf;
			{9'd282, 8'd133}: color_data = 12'h0be;
			{9'd282, 8'd134}: color_data = 12'h056;
			{9'd282, 8'd135}: color_data = 12'h012;
			{9'd282, 8'd136}: color_data = 12'h08b;
			{9'd282, 8'd137}: color_data = 12'h034;
			{9'd282, 8'd170}: color_data = 12'h000;
			{9'd282, 8'd171}: color_data = 12'h068;
			{9'd282, 8'd172}: color_data = 12'h8ef;
			{9'd282, 8'd173}: color_data = 12'hdff;
			{9'd282, 8'd174}: color_data = 12'h4cf;
			{9'd282, 8'd175}: color_data = 12'h0cf;
			{9'd282, 8'd176}: color_data = 12'h0ae;
			{9'd282, 8'd177}: color_data = 12'h035;
			{9'd282, 8'd178}: color_data = 12'h023;
			{9'd282, 8'd179}: color_data = 12'h08c;
			{9'd282, 8'd180}: color_data = 12'h023;
			{9'd282, 8'd222}: color_data = 12'h200;
			{9'd282, 8'd223}: color_data = 12'h900;
			{9'd282, 8'd224}: color_data = 12'hb00;
			{9'd282, 8'd225}: color_data = 12'h800;
			{9'd282, 8'd226}: color_data = 12'h200;
			{9'd282, 8'd227}: color_data = 12'hb30;
			{9'd282, 8'd228}: color_data = 12'hc10;
			{9'd282, 8'd229}: color_data = 12'h800;
			{9'd282, 8'd230}: color_data = 12'h300;
			{9'd282, 8'd231}: color_data = 12'h400;
			{9'd282, 8'd232}: color_data = 12'ha00;
			{9'd282, 8'd233}: color_data = 12'ha00;
			{9'd282, 8'd234}: color_data = 12'h500;
			{9'd282, 8'd235}: color_data = 12'h510;
			{9'd282, 8'd236}: color_data = 12'hd30;
			{9'd282, 8'd237}: color_data = 12'ha00;
			{9'd282, 8'd238}: color_data = 12'h700;
			{9'd282, 8'd239}: color_data = 12'h100;
			{9'd283, 8'd15}: color_data = 12'h110;
			{9'd283, 8'd16}: color_data = 12'h890;
			{9'd283, 8'd17}: color_data = 12'had1;
			{9'd283, 8'd18}: color_data = 12'hefb;
			{9'd283, 8'd19}: color_data = 12'hfff;
			{9'd283, 8'd20}: color_data = 12'hcd6;
			{9'd283, 8'd21}: color_data = 12'h9b0;
			{9'd283, 8'd22}: color_data = 12'hac0;
			{9'd283, 8'd23}: color_data = 12'hac0;
			{9'd283, 8'd24}: color_data = 12'hac0;
			{9'd283, 8'd25}: color_data = 12'hac0;
			{9'd283, 8'd26}: color_data = 12'h9b0;
			{9'd283, 8'd27}: color_data = 12'h550;
			{9'd283, 8'd28}: color_data = 12'h020;
			{9'd283, 8'd29}: color_data = 12'h140;
			{9'd283, 8'd30}: color_data = 12'h240;
			{9'd283, 8'd31}: color_data = 12'h660;
			{9'd283, 8'd32}: color_data = 12'h760;
			{9'd283, 8'd33}: color_data = 12'h120;
			{9'd283, 8'd68}: color_data = 12'h047;
			{9'd283, 8'd69}: color_data = 12'h6df;
			{9'd283, 8'd70}: color_data = 12'hfff;
			{9'd283, 8'd71}: color_data = 12'hdff;
			{9'd283, 8'd72}: color_data = 12'h5df;
			{9'd283, 8'd73}: color_data = 12'h068;
			{9'd283, 8'd74}: color_data = 12'h000;
			{9'd283, 8'd75}: color_data = 12'h012;
			{9'd283, 8'd76}: color_data = 12'h08c;
			{9'd283, 8'd77}: color_data = 12'h034;
			{9'd283, 8'd128}: color_data = 12'h047;
			{9'd283, 8'd129}: color_data = 12'h6df;
			{9'd283, 8'd130}: color_data = 12'hfff;
			{9'd283, 8'd131}: color_data = 12'hdff;
			{9'd283, 8'd132}: color_data = 12'h5df;
			{9'd283, 8'd133}: color_data = 12'h068;
			{9'd283, 8'd134}: color_data = 12'h000;
			{9'd283, 8'd135}: color_data = 12'h012;
			{9'd283, 8'd136}: color_data = 12'h08c;
			{9'd283, 8'd137}: color_data = 12'h034;
			{9'd283, 8'd170}: color_data = 12'h000;
			{9'd283, 8'd171}: color_data = 12'h068;
			{9'd283, 8'd172}: color_data = 12'h8ef;
			{9'd283, 8'd173}: color_data = 12'hfff;
			{9'd283, 8'd174}: color_data = 12'hcff;
			{9'd283, 8'd175}: color_data = 12'h4ce;
			{9'd283, 8'd176}: color_data = 12'h057;
			{9'd283, 8'd177}: color_data = 12'h000;
			{9'd283, 8'd178}: color_data = 12'h023;
			{9'd283, 8'd179}: color_data = 12'h08c;
			{9'd283, 8'd180}: color_data = 12'h023;
			{9'd283, 8'd222}: color_data = 12'h200;
			{9'd283, 8'd223}: color_data = 12'h900;
			{9'd283, 8'd224}: color_data = 12'ha00;
			{9'd283, 8'd225}: color_data = 12'h700;
			{9'd283, 8'd226}: color_data = 12'h200;
			{9'd283, 8'd227}: color_data = 12'hb30;
			{9'd283, 8'd228}: color_data = 12'he20;
			{9'd283, 8'd229}: color_data = 12'ha00;
			{9'd283, 8'd230}: color_data = 12'h300;
			{9'd283, 8'd231}: color_data = 12'h400;
			{9'd283, 8'd232}: color_data = 12'ha00;
			{9'd283, 8'd233}: color_data = 12'ha00;
			{9'd283, 8'd234}: color_data = 12'h400;
			{9'd283, 8'd235}: color_data = 12'h510;
			{9'd283, 8'd236}: color_data = 12'hf40;
			{9'd283, 8'd237}: color_data = 12'hd10;
			{9'd283, 8'd238}: color_data = 12'h800;
			{9'd283, 8'd239}: color_data = 12'h100;
			{9'd284, 8'd15}: color_data = 12'h010;
			{9'd284, 8'd16}: color_data = 12'h670;
			{9'd284, 8'd17}: color_data = 12'h8a0;
			{9'd284, 8'd18}: color_data = 12'hbc9;
			{9'd284, 8'd19}: color_data = 12'hcdd;
			{9'd284, 8'd20}: color_data = 12'h9a4;
			{9'd284, 8'd21}: color_data = 12'h690;
			{9'd284, 8'd22}: color_data = 12'h790;
			{9'd284, 8'd23}: color_data = 12'h790;
			{9'd284, 8'd24}: color_data = 12'h790;
			{9'd284, 8'd25}: color_data = 12'h7a0;
			{9'd284, 8'd26}: color_data = 12'h780;
			{9'd284, 8'd27}: color_data = 12'h440;
			{9'd284, 8'd28}: color_data = 12'h020;
			{9'd284, 8'd29}: color_data = 12'h130;
			{9'd284, 8'd30}: color_data = 12'h140;
			{9'd284, 8'd31}: color_data = 12'h450;
			{9'd284, 8'd32}: color_data = 12'h550;
			{9'd284, 8'd33}: color_data = 12'h110;
			{9'd284, 8'd68}: color_data = 12'h047;
			{9'd284, 8'd69}: color_data = 12'h6df;
			{9'd284, 8'd70}: color_data = 12'hfff;
			{9'd284, 8'd71}: color_data = 12'hfff;
			{9'd284, 8'd72}: color_data = 12'h9aa;
			{9'd284, 8'd73}: color_data = 12'h011;
			{9'd284, 8'd75}: color_data = 12'h012;
			{9'd284, 8'd76}: color_data = 12'h08c;
			{9'd284, 8'd77}: color_data = 12'h034;
			{9'd284, 8'd128}: color_data = 12'h047;
			{9'd284, 8'd129}: color_data = 12'h6df;
			{9'd284, 8'd130}: color_data = 12'hfff;
			{9'd284, 8'd131}: color_data = 12'hfff;
			{9'd284, 8'd132}: color_data = 12'h9aa;
			{9'd284, 8'd133}: color_data = 12'h111;
			{9'd284, 8'd135}: color_data = 12'h012;
			{9'd284, 8'd136}: color_data = 12'h08c;
			{9'd284, 8'd137}: color_data = 12'h034;
			{9'd284, 8'd170}: color_data = 12'h000;
			{9'd284, 8'd171}: color_data = 12'h068;
			{9'd284, 8'd172}: color_data = 12'h7ef;
			{9'd284, 8'd173}: color_data = 12'hfff;
			{9'd284, 8'd174}: color_data = 12'hfff;
			{9'd284, 8'd175}: color_data = 12'h899;
			{9'd284, 8'd176}: color_data = 12'h001;
			{9'd284, 8'd178}: color_data = 12'h024;
			{9'd284, 8'd179}: color_data = 12'h08c;
			{9'd284, 8'd180}: color_data = 12'h023;
			{9'd284, 8'd222}: color_data = 12'h200;
			{9'd284, 8'd223}: color_data = 12'h800;
			{9'd284, 8'd224}: color_data = 12'ha00;
			{9'd284, 8'd225}: color_data = 12'h800;
			{9'd284, 8'd226}: color_data = 12'h200;
			{9'd284, 8'd227}: color_data = 12'h930;
			{9'd284, 8'd228}: color_data = 12'hd30;
			{9'd284, 8'd229}: color_data = 12'h910;
			{9'd284, 8'd230}: color_data = 12'h200;
			{9'd284, 8'd231}: color_data = 12'h400;
			{9'd284, 8'd232}: color_data = 12'h900;
			{9'd284, 8'd233}: color_data = 12'ha00;
			{9'd284, 8'd234}: color_data = 12'h400;
			{9'd284, 8'd235}: color_data = 12'h310;
			{9'd284, 8'd236}: color_data = 12'hc30;
			{9'd284, 8'd237}: color_data = 12'hc20;
			{9'd284, 8'd238}: color_data = 12'h600;
			{9'd284, 8'd239}: color_data = 12'h000;
			{9'd285, 8'd15}: color_data = 12'h000;
			{9'd285, 8'd16}: color_data = 12'h110;
			{9'd285, 8'd17}: color_data = 12'h130;
			{9'd285, 8'd18}: color_data = 12'h242;
			{9'd285, 8'd19}: color_data = 12'h343;
			{9'd285, 8'd20}: color_data = 12'h242;
			{9'd285, 8'd21}: color_data = 12'h130;
			{9'd285, 8'd22}: color_data = 12'h130;
			{9'd285, 8'd23}: color_data = 12'h130;
			{9'd285, 8'd24}: color_data = 12'h130;
			{9'd285, 8'd25}: color_data = 12'h130;
			{9'd285, 8'd26}: color_data = 12'h130;
			{9'd285, 8'd27}: color_data = 12'h020;
			{9'd285, 8'd28}: color_data = 12'h020;
			{9'd285, 8'd29}: color_data = 12'h020;
			{9'd285, 8'd30}: color_data = 12'h020;
			{9'd285, 8'd31}: color_data = 12'h120;
			{9'd285, 8'd32}: color_data = 12'h110;
			{9'd285, 8'd33}: color_data = 12'h000;
			{9'd285, 8'd68}: color_data = 12'h047;
			{9'd285, 8'd69}: color_data = 12'h6df;
			{9'd285, 8'd70}: color_data = 12'hfff;
			{9'd285, 8'd71}: color_data = 12'hcbb;
			{9'd285, 8'd72}: color_data = 12'h323;
			{9'd285, 8'd73}: color_data = 12'h002;
			{9'd285, 8'd74}: color_data = 12'h000;
			{9'd285, 8'd75}: color_data = 12'h012;
			{9'd285, 8'd76}: color_data = 12'h08c;
			{9'd285, 8'd77}: color_data = 12'h034;
			{9'd285, 8'd128}: color_data = 12'h047;
			{9'd285, 8'd129}: color_data = 12'h6df;
			{9'd285, 8'd130}: color_data = 12'hfff;
			{9'd285, 8'd131}: color_data = 12'hcbb;
			{9'd285, 8'd132}: color_data = 12'h323;
			{9'd285, 8'd133}: color_data = 12'h002;
			{9'd285, 8'd134}: color_data = 12'h000;
			{9'd285, 8'd135}: color_data = 12'h012;
			{9'd285, 8'd136}: color_data = 12'h08c;
			{9'd285, 8'd137}: color_data = 12'h034;
			{9'd285, 8'd170}: color_data = 12'h000;
			{9'd285, 8'd171}: color_data = 12'h068;
			{9'd285, 8'd172}: color_data = 12'h8ef;
			{9'd285, 8'd173}: color_data = 12'hfff;
			{9'd285, 8'd174}: color_data = 12'haa9;
			{9'd285, 8'd175}: color_data = 12'h212;
			{9'd285, 8'd176}: color_data = 12'h002;
			{9'd285, 8'd178}: color_data = 12'h023;
			{9'd285, 8'd179}: color_data = 12'h08c;
			{9'd285, 8'd180}: color_data = 12'h023;
			{9'd285, 8'd222}: color_data = 12'h200;
			{9'd285, 8'd223}: color_data = 12'h900;
			{9'd285, 8'd224}: color_data = 12'ha00;
			{9'd285, 8'd225}: color_data = 12'h800;
			{9'd285, 8'd226}: color_data = 12'h100;
			{9'd285, 8'd227}: color_data = 12'h100;
			{9'd285, 8'd228}: color_data = 12'h300;
			{9'd285, 8'd229}: color_data = 12'h200;
			{9'd285, 8'd230}: color_data = 12'h000;
			{9'd285, 8'd231}: color_data = 12'h500;
			{9'd285, 8'd232}: color_data = 12'ha00;
			{9'd285, 8'd233}: color_data = 12'ha00;
			{9'd285, 8'd234}: color_data = 12'h500;
			{9'd285, 8'd235}: color_data = 12'h000;
			{9'd285, 8'd236}: color_data = 12'h200;
			{9'd285, 8'd237}: color_data = 12'h300;
			{9'd285, 8'd238}: color_data = 12'h100;
			{9'd285, 8'd239}: color_data = 12'h000;
			{9'd286, 8'd16}: color_data = 12'h000;
			{9'd286, 8'd17}: color_data = 12'h230;
			{9'd286, 8'd18}: color_data = 12'h340;
			{9'd286, 8'd19}: color_data = 12'h786;
			{9'd286, 8'd20}: color_data = 12'habb;
			{9'd286, 8'd21}: color_data = 12'h674;
			{9'd286, 8'd22}: color_data = 12'h330;
			{9'd286, 8'd23}: color_data = 12'h340;
			{9'd286, 8'd24}: color_data = 12'h340;
			{9'd286, 8'd25}: color_data = 12'h440;
			{9'd286, 8'd26}: color_data = 12'h230;
			{9'd286, 8'd27}: color_data = 12'h020;
			{9'd286, 8'd28}: color_data = 12'h030;
			{9'd286, 8'd29}: color_data = 12'h130;
			{9'd286, 8'd30}: color_data = 12'h440;
			{9'd286, 8'd31}: color_data = 12'h440;
			{9'd286, 8'd32}: color_data = 12'h010;
			{9'd286, 8'd68}: color_data = 12'h047;
			{9'd286, 8'd69}: color_data = 12'h6ef;
			{9'd286, 8'd70}: color_data = 12'hccc;
			{9'd286, 8'd71}: color_data = 12'h434;
			{9'd286, 8'd72}: color_data = 12'h003;
			{9'd286, 8'd73}: color_data = 12'h005;
			{9'd286, 8'd74}: color_data = 12'h002;
			{9'd286, 8'd75}: color_data = 12'h012;
			{9'd286, 8'd76}: color_data = 12'h08c;
			{9'd286, 8'd77}: color_data = 12'h034;
			{9'd286, 8'd128}: color_data = 12'h047;
			{9'd286, 8'd129}: color_data = 12'h6ef;
			{9'd286, 8'd130}: color_data = 12'hddc;
			{9'd286, 8'd131}: color_data = 12'h434;
			{9'd286, 8'd132}: color_data = 12'h003;
			{9'd286, 8'd133}: color_data = 12'h005;
			{9'd286, 8'd134}: color_data = 12'h002;
			{9'd286, 8'd135}: color_data = 12'h012;
			{9'd286, 8'd136}: color_data = 12'h08c;
			{9'd286, 8'd137}: color_data = 12'h034;
			{9'd286, 8'd170}: color_data = 12'h000;
			{9'd286, 8'd171}: color_data = 12'h068;
			{9'd286, 8'd172}: color_data = 12'h8ff;
			{9'd286, 8'd173}: color_data = 12'hcbb;
			{9'd286, 8'd174}: color_data = 12'h223;
			{9'd286, 8'd175}: color_data = 12'h003;
			{9'd286, 8'd176}: color_data = 12'h005;
			{9'd286, 8'd177}: color_data = 12'h002;
			{9'd286, 8'd178}: color_data = 12'h023;
			{9'd286, 8'd179}: color_data = 12'h09c;
			{9'd286, 8'd180}: color_data = 12'h023;
			{9'd286, 8'd222}: color_data = 12'h300;
			{9'd286, 8'd223}: color_data = 12'hc20;
			{9'd286, 8'd224}: color_data = 12'ha00;
			{9'd286, 8'd225}: color_data = 12'h800;
			{9'd286, 8'd226}: color_data = 12'h100;
			{9'd286, 8'd227}: color_data = 12'h300;
			{9'd286, 8'd228}: color_data = 12'h500;
			{9'd286, 8'd229}: color_data = 12'h500;
			{9'd286, 8'd230}: color_data = 12'h100;
			{9'd286, 8'd231}: color_data = 12'h710;
			{9'd286, 8'd232}: color_data = 12'hc10;
			{9'd286, 8'd233}: color_data = 12'h900;
			{9'd286, 8'd234}: color_data = 12'h500;
			{9'd286, 8'd235}: color_data = 12'h100;
			{9'd286, 8'd236}: color_data = 12'h500;
			{9'd286, 8'd237}: color_data = 12'h600;
			{9'd286, 8'd238}: color_data = 12'h400;
			{9'd286, 8'd239}: color_data = 12'h000;
			{9'd287, 8'd16}: color_data = 12'h000;
			{9'd287, 8'd17}: color_data = 12'h670;
			{9'd287, 8'd18}: color_data = 12'h890;
			{9'd287, 8'd19}: color_data = 12'hdda;
			{9'd287, 8'd20}: color_data = 12'hfff;
			{9'd287, 8'd21}: color_data = 12'hbc7;
			{9'd287, 8'd22}: color_data = 12'h780;
			{9'd287, 8'd23}: color_data = 12'h890;
			{9'd287, 8'd24}: color_data = 12'h890;
			{9'd287, 8'd25}: color_data = 12'h880;
			{9'd287, 8'd26}: color_data = 12'h450;
			{9'd287, 8'd27}: color_data = 12'h020;
			{9'd287, 8'd28}: color_data = 12'h140;
			{9'd287, 8'd29}: color_data = 12'h250;
			{9'd287, 8'd30}: color_data = 12'h660;
			{9'd287, 8'd31}: color_data = 12'h660;
			{9'd287, 8'd32}: color_data = 12'h110;
			{9'd287, 8'd68}: color_data = 12'h057;
			{9'd287, 8'd69}: color_data = 12'h3bd;
			{9'd287, 8'd70}: color_data = 12'h555;
			{9'd287, 8'd71}: color_data = 12'h002;
			{9'd287, 8'd72}: color_data = 12'h005;
			{9'd287, 8'd73}: color_data = 12'h005;
			{9'd287, 8'd74}: color_data = 12'h004;
			{9'd287, 8'd75}: color_data = 12'h025;
			{9'd287, 8'd76}: color_data = 12'h09c;
			{9'd287, 8'd77}: color_data = 12'h034;
			{9'd287, 8'd128}: color_data = 12'h057;
			{9'd287, 8'd129}: color_data = 12'h3bd;
			{9'd287, 8'd130}: color_data = 12'h555;
			{9'd287, 8'd131}: color_data = 12'h002;
			{9'd287, 8'd132}: color_data = 12'h005;
			{9'd287, 8'd133}: color_data = 12'h005;
			{9'd287, 8'd134}: color_data = 12'h004;
			{9'd287, 8'd135}: color_data = 12'h025;
			{9'd287, 8'd136}: color_data = 12'h09c;
			{9'd287, 8'd137}: color_data = 12'h034;
			{9'd287, 8'd170}: color_data = 12'h000;
			{9'd287, 8'd171}: color_data = 12'h079;
			{9'd287, 8'd172}: color_data = 12'h4bd;
			{9'd287, 8'd173}: color_data = 12'h444;
			{9'd287, 8'd174}: color_data = 12'h002;
			{9'd287, 8'd175}: color_data = 12'h005;
			{9'd287, 8'd176}: color_data = 12'h005;
			{9'd287, 8'd177}: color_data = 12'h004;
			{9'd287, 8'd178}: color_data = 12'h036;
			{9'd287, 8'd179}: color_data = 12'h09c;
			{9'd287, 8'd180}: color_data = 12'h023;
			{9'd287, 8'd222}: color_data = 12'h410;
			{9'd287, 8'd223}: color_data = 12'hd30;
			{9'd287, 8'd224}: color_data = 12'hb00;
			{9'd287, 8'd225}: color_data = 12'h700;
			{9'd287, 8'd226}: color_data = 12'h200;
			{9'd287, 8'd227}: color_data = 12'h700;
			{9'd287, 8'd228}: color_data = 12'hb00;
			{9'd287, 8'd229}: color_data = 12'ha00;
			{9'd287, 8'd230}: color_data = 12'h300;
			{9'd287, 8'd231}: color_data = 12'h820;
			{9'd287, 8'd232}: color_data = 12'hd20;
			{9'd287, 8'd233}: color_data = 12'h900;
			{9'd287, 8'd234}: color_data = 12'h500;
			{9'd287, 8'd235}: color_data = 12'h300;
			{9'd287, 8'd236}: color_data = 12'h900;
			{9'd287, 8'd237}: color_data = 12'hb00;
			{9'd287, 8'd238}: color_data = 12'h800;
			{9'd287, 8'd239}: color_data = 12'h100;
			{9'd288, 8'd16}: color_data = 12'h010;
			{9'd288, 8'd17}: color_data = 12'h780;
			{9'd288, 8'd18}: color_data = 12'hac0;
			{9'd288, 8'd19}: color_data = 12'hdea;
			{9'd288, 8'd20}: color_data = 12'hfff;
			{9'd288, 8'd21}: color_data = 12'hcd7;
			{9'd288, 8'd22}: color_data = 12'h9b0;
			{9'd288, 8'd23}: color_data = 12'h9b0;
			{9'd288, 8'd24}: color_data = 12'h9c0;
			{9'd288, 8'd25}: color_data = 12'h9a0;
			{9'd288, 8'd26}: color_data = 12'h450;
			{9'd288, 8'd27}: color_data = 12'h020;
			{9'd288, 8'd28}: color_data = 12'h140;
			{9'd288, 8'd29}: color_data = 12'h240;
			{9'd288, 8'd30}: color_data = 12'h660;
			{9'd288, 8'd31}: color_data = 12'h660;
			{9'd288, 8'd32}: color_data = 12'h110;
			{9'd288, 8'd68}: color_data = 12'h035;
			{9'd288, 8'd69}: color_data = 12'h047;
			{9'd288, 8'd70}: color_data = 12'h001;
			{9'd288, 8'd71}: color_data = 12'h004;
			{9'd288, 8'd72}: color_data = 12'h004;
			{9'd288, 8'd73}: color_data = 12'h004;
			{9'd288, 8'd74}: color_data = 12'h004;
			{9'd288, 8'd75}: color_data = 12'h015;
			{9'd288, 8'd76}: color_data = 12'h059;
			{9'd288, 8'd77}: color_data = 12'h023;
			{9'd288, 8'd128}: color_data = 12'h035;
			{9'd288, 8'd129}: color_data = 12'h047;
			{9'd288, 8'd130}: color_data = 12'h001;
			{9'd288, 8'd131}: color_data = 12'h004;
			{9'd288, 8'd132}: color_data = 12'h004;
			{9'd288, 8'd133}: color_data = 12'h004;
			{9'd288, 8'd134}: color_data = 12'h004;
			{9'd288, 8'd135}: color_data = 12'h015;
			{9'd288, 8'd136}: color_data = 12'h059;
			{9'd288, 8'd137}: color_data = 12'h023;
			{9'd288, 8'd170}: color_data = 12'h000;
			{9'd288, 8'd171}: color_data = 12'h047;
			{9'd288, 8'd172}: color_data = 12'h036;
			{9'd288, 8'd173}: color_data = 12'h001;
			{9'd288, 8'd174}: color_data = 12'h004;
			{9'd288, 8'd175}: color_data = 12'h004;
			{9'd288, 8'd176}: color_data = 12'h004;
			{9'd288, 8'd177}: color_data = 12'h004;
			{9'd288, 8'd178}: color_data = 12'h016;
			{9'd288, 8'd179}: color_data = 12'h059;
			{9'd288, 8'd180}: color_data = 12'h012;
			{9'd288, 8'd222}: color_data = 12'h410;
			{9'd288, 8'd223}: color_data = 12'he40;
			{9'd288, 8'd224}: color_data = 12'hd20;
			{9'd288, 8'd225}: color_data = 12'h800;
			{9'd288, 8'd226}: color_data = 12'h200;
			{9'd288, 8'd227}: color_data = 12'h600;
			{9'd288, 8'd228}: color_data = 12'ha00;
			{9'd288, 8'd229}: color_data = 12'h900;
			{9'd288, 8'd230}: color_data = 12'h300;
			{9'd288, 8'd231}: color_data = 12'h820;
			{9'd288, 8'd232}: color_data = 12'hf30;
			{9'd288, 8'd233}: color_data = 12'hc00;
			{9'd288, 8'd234}: color_data = 12'h500;
			{9'd288, 8'd235}: color_data = 12'h200;
			{9'd288, 8'd236}: color_data = 12'h900;
			{9'd288, 8'd237}: color_data = 12'ha00;
			{9'd288, 8'd238}: color_data = 12'h700;
			{9'd288, 8'd239}: color_data = 12'h100;
			{9'd289, 8'd16}: color_data = 12'h010;
			{9'd289, 8'd17}: color_data = 12'h780;
			{9'd289, 8'd18}: color_data = 12'hac0;
			{9'd289, 8'd19}: color_data = 12'hdea;
			{9'd289, 8'd20}: color_data = 12'hfff;
			{9'd289, 8'd21}: color_data = 12'hcd7;
			{9'd289, 8'd22}: color_data = 12'h9b0;
			{9'd289, 8'd23}: color_data = 12'h9b0;
			{9'd289, 8'd24}: color_data = 12'h9c0;
			{9'd289, 8'd25}: color_data = 12'h8a0;
			{9'd289, 8'd26}: color_data = 12'h450;
			{9'd289, 8'd27}: color_data = 12'h020;
			{9'd289, 8'd28}: color_data = 12'h140;
			{9'd289, 8'd29}: color_data = 12'h240;
			{9'd289, 8'd30}: color_data = 12'h660;
			{9'd289, 8'd31}: color_data = 12'h660;
			{9'd289, 8'd32}: color_data = 12'h110;
			{9'd289, 8'd68}: color_data = 12'h013;
			{9'd289, 8'd69}: color_data = 12'h027;
			{9'd289, 8'd70}: color_data = 12'h016;
			{9'd289, 8'd71}: color_data = 12'h027;
			{9'd289, 8'd72}: color_data = 12'h027;
			{9'd289, 8'd73}: color_data = 12'h027;
			{9'd289, 8'd74}: color_data = 12'h027;
			{9'd289, 8'd75}: color_data = 12'h028;
			{9'd289, 8'd76}: color_data = 12'h027;
			{9'd289, 8'd77}: color_data = 12'h001;
			{9'd289, 8'd128}: color_data = 12'h013;
			{9'd289, 8'd129}: color_data = 12'h027;
			{9'd289, 8'd130}: color_data = 12'h016;
			{9'd289, 8'd131}: color_data = 12'h027;
			{9'd289, 8'd132}: color_data = 12'h027;
			{9'd289, 8'd133}: color_data = 12'h017;
			{9'd289, 8'd134}: color_data = 12'h027;
			{9'd289, 8'd135}: color_data = 12'h028;
			{9'd289, 8'd136}: color_data = 12'h027;
			{9'd289, 8'd137}: color_data = 12'h001;
			{9'd289, 8'd170}: color_data = 12'h000;
			{9'd289, 8'd171}: color_data = 12'h014;
			{9'd289, 8'd172}: color_data = 12'h027;
			{9'd289, 8'd173}: color_data = 12'h016;
			{9'd289, 8'd174}: color_data = 12'h027;
			{9'd289, 8'd175}: color_data = 12'h027;
			{9'd289, 8'd176}: color_data = 12'h027;
			{9'd289, 8'd177}: color_data = 12'h027;
			{9'd289, 8'd178}: color_data = 12'h028;
			{9'd289, 8'd179}: color_data = 12'h026;
			{9'd289, 8'd180}: color_data = 12'h001;
			{9'd289, 8'd222}: color_data = 12'h300;
			{9'd289, 8'd223}: color_data = 12'hc30;
			{9'd289, 8'd224}: color_data = 12'hc30;
			{9'd289, 8'd225}: color_data = 12'h600;
			{9'd289, 8'd226}: color_data = 12'h100;
			{9'd289, 8'd227}: color_data = 12'h600;
			{9'd289, 8'd228}: color_data = 12'ha00;
			{9'd289, 8'd229}: color_data = 12'h900;
			{9'd289, 8'd230}: color_data = 12'h300;
			{9'd289, 8'd231}: color_data = 12'h620;
			{9'd289, 8'd232}: color_data = 12'hd40;
			{9'd289, 8'd233}: color_data = 12'ha20;
			{9'd289, 8'd234}: color_data = 12'h300;
			{9'd289, 8'd235}: color_data = 12'h200;
			{9'd289, 8'd236}: color_data = 12'h900;
			{9'd289, 8'd237}: color_data = 12'ha00;
			{9'd289, 8'd238}: color_data = 12'h700;
			{9'd289, 8'd239}: color_data = 12'h100;
			{9'd290, 8'd16}: color_data = 12'h010;
			{9'd290, 8'd17}: color_data = 12'h780;
			{9'd290, 8'd18}: color_data = 12'hac0;
			{9'd290, 8'd19}: color_data = 12'hdea;
			{9'd290, 8'd20}: color_data = 12'hfff;
			{9'd290, 8'd21}: color_data = 12'hcd7;
			{9'd290, 8'd22}: color_data = 12'h9b0;
			{9'd290, 8'd23}: color_data = 12'h9b0;
			{9'd290, 8'd24}: color_data = 12'h9b0;
			{9'd290, 8'd25}: color_data = 12'h8a0;
			{9'd290, 8'd26}: color_data = 12'h450;
			{9'd290, 8'd27}: color_data = 12'h020;
			{9'd290, 8'd28}: color_data = 12'h140;
			{9'd290, 8'd29}: color_data = 12'h240;
			{9'd290, 8'd30}: color_data = 12'h660;
			{9'd290, 8'd31}: color_data = 12'h660;
			{9'd290, 8'd32}: color_data = 12'h110;
			{9'd290, 8'd68}: color_data = 12'h036;
			{9'd290, 8'd69}: color_data = 12'h09e;
			{9'd290, 8'd70}: color_data = 12'h09e;
			{9'd290, 8'd71}: color_data = 12'h09e;
			{9'd290, 8'd72}: color_data = 12'h09e;
			{9'd290, 8'd73}: color_data = 12'h09e;
			{9'd290, 8'd74}: color_data = 12'h09e;
			{9'd290, 8'd75}: color_data = 12'h09e;
			{9'd290, 8'd76}: color_data = 12'h08c;
			{9'd290, 8'd77}: color_data = 12'h023;
			{9'd290, 8'd128}: color_data = 12'h035;
			{9'd290, 8'd129}: color_data = 12'h09e;
			{9'd290, 8'd130}: color_data = 12'h09e;
			{9'd290, 8'd131}: color_data = 12'h09e;
			{9'd290, 8'd132}: color_data = 12'h09e;
			{9'd290, 8'd133}: color_data = 12'h09e;
			{9'd290, 8'd134}: color_data = 12'h09e;
			{9'd290, 8'd135}: color_data = 12'h09e;
			{9'd290, 8'd136}: color_data = 12'h08c;
			{9'd290, 8'd137}: color_data = 12'h023;
			{9'd290, 8'd170}: color_data = 12'h000;
			{9'd290, 8'd171}: color_data = 12'h057;
			{9'd290, 8'd172}: color_data = 12'h0ae;
			{9'd290, 8'd173}: color_data = 12'h09e;
			{9'd290, 8'd174}: color_data = 12'h09e;
			{9'd290, 8'd175}: color_data = 12'h09e;
			{9'd290, 8'd176}: color_data = 12'h09e;
			{9'd290, 8'd177}: color_data = 12'h09e;
			{9'd290, 8'd178}: color_data = 12'h09e;
			{9'd290, 8'd179}: color_data = 12'h07b;
			{9'd290, 8'd180}: color_data = 12'h012;
			{9'd290, 8'd222}: color_data = 12'h000;
			{9'd290, 8'd223}: color_data = 12'h200;
			{9'd290, 8'd224}: color_data = 12'h300;
			{9'd290, 8'd225}: color_data = 12'h100;
			{9'd290, 8'd226}: color_data = 12'h000;
			{9'd290, 8'd227}: color_data = 12'h700;
			{9'd290, 8'd228}: color_data = 12'ha00;
			{9'd290, 8'd229}: color_data = 12'h900;
			{9'd290, 8'd230}: color_data = 12'h300;
			{9'd290, 8'd231}: color_data = 12'h100;
			{9'd290, 8'd232}: color_data = 12'h310;
			{9'd290, 8'd233}: color_data = 12'h200;
			{9'd290, 8'd234}: color_data = 12'h000;
			{9'd290, 8'd235}: color_data = 12'h300;
			{9'd290, 8'd236}: color_data = 12'h900;
			{9'd290, 8'd237}: color_data = 12'ha00;
			{9'd290, 8'd238}: color_data = 12'h700;
			{9'd290, 8'd239}: color_data = 12'h100;
			{9'd291, 8'd16}: color_data = 12'h010;
			{9'd291, 8'd17}: color_data = 12'h780;
			{9'd291, 8'd18}: color_data = 12'hac0;
			{9'd291, 8'd19}: color_data = 12'hdea;
			{9'd291, 8'd20}: color_data = 12'hfff;
			{9'd291, 8'd21}: color_data = 12'hcd7;
			{9'd291, 8'd22}: color_data = 12'h9b0;
			{9'd291, 8'd23}: color_data = 12'h9b0;
			{9'd291, 8'd24}: color_data = 12'h9b0;
			{9'd291, 8'd25}: color_data = 12'h8a0;
			{9'd291, 8'd26}: color_data = 12'h450;
			{9'd291, 8'd27}: color_data = 12'h020;
			{9'd291, 8'd28}: color_data = 12'h140;
			{9'd291, 8'd29}: color_data = 12'h240;
			{9'd291, 8'd30}: color_data = 12'h660;
			{9'd291, 8'd31}: color_data = 12'h660;
			{9'd291, 8'd32}: color_data = 12'h110;
			{9'd291, 8'd68}: color_data = 12'h057;
			{9'd291, 8'd69}: color_data = 12'h4ef;
			{9'd291, 8'd70}: color_data = 12'h7ef;
			{9'd291, 8'd71}: color_data = 12'h0cf;
			{9'd291, 8'd72}: color_data = 12'h0cf;
			{9'd291, 8'd73}: color_data = 12'h0df;
			{9'd291, 8'd74}: color_data = 12'h0bd;
			{9'd291, 8'd75}: color_data = 12'h068;
			{9'd291, 8'd76}: color_data = 12'h09c;
			{9'd291, 8'd77}: color_data = 12'h034;
			{9'd291, 8'd128}: color_data = 12'h057;
			{9'd291, 8'd129}: color_data = 12'h4ef;
			{9'd291, 8'd130}: color_data = 12'h7ef;
			{9'd291, 8'd131}: color_data = 12'h0cf;
			{9'd291, 8'd132}: color_data = 12'h0cf;
			{9'd291, 8'd133}: color_data = 12'h0df;
			{9'd291, 8'd134}: color_data = 12'h0bd;
			{9'd291, 8'd135}: color_data = 12'h068;
			{9'd291, 8'd136}: color_data = 12'h09c;
			{9'd291, 8'd137}: color_data = 12'h034;
			{9'd291, 8'd170}: color_data = 12'h000;
			{9'd291, 8'd171}: color_data = 12'h069;
			{9'd291, 8'd172}: color_data = 12'h6ef;
			{9'd291, 8'd173}: color_data = 12'h6ef;
			{9'd291, 8'd174}: color_data = 12'h0cf;
			{9'd291, 8'd175}: color_data = 12'h0cf;
			{9'd291, 8'd176}: color_data = 12'h0df;
			{9'd291, 8'd177}: color_data = 12'h0ac;
			{9'd291, 8'd178}: color_data = 12'h079;
			{9'd291, 8'd179}: color_data = 12'h09c;
			{9'd291, 8'd180}: color_data = 12'h023;
			{9'd291, 8'd222}: color_data = 12'h100;
			{9'd291, 8'd223}: color_data = 12'h500;
			{9'd291, 8'd224}: color_data = 12'h500;
			{9'd291, 8'd225}: color_data = 12'h400;
			{9'd291, 8'd226}: color_data = 12'h200;
			{9'd291, 8'd227}: color_data = 12'ha20;
			{9'd291, 8'd228}: color_data = 12'hb10;
			{9'd291, 8'd229}: color_data = 12'h900;
			{9'd291, 8'd230}: color_data = 12'h300;
			{9'd291, 8'd231}: color_data = 12'h200;
			{9'd291, 8'd232}: color_data = 12'h500;
			{9'd291, 8'd233}: color_data = 12'h500;
			{9'd291, 8'd234}: color_data = 12'h200;
			{9'd291, 8'd235}: color_data = 12'h410;
			{9'd291, 8'd236}: color_data = 12'hc20;
			{9'd291, 8'd237}: color_data = 12'ha00;
			{9'd291, 8'd238}: color_data = 12'h700;
			{9'd291, 8'd239}: color_data = 12'h100;
			{9'd292, 8'd16}: color_data = 12'h010;
			{9'd292, 8'd17}: color_data = 12'h780;
			{9'd292, 8'd18}: color_data = 12'hac0;
			{9'd292, 8'd19}: color_data = 12'hdea;
			{9'd292, 8'd20}: color_data = 12'hfff;
			{9'd292, 8'd21}: color_data = 12'hcd7;
			{9'd292, 8'd22}: color_data = 12'h9b0;
			{9'd292, 8'd23}: color_data = 12'h9b0;
			{9'd292, 8'd24}: color_data = 12'h9b0;
			{9'd292, 8'd25}: color_data = 12'h8a0;
			{9'd292, 8'd26}: color_data = 12'h450;
			{9'd292, 8'd27}: color_data = 12'h020;
			{9'd292, 8'd28}: color_data = 12'h140;
			{9'd292, 8'd29}: color_data = 12'h240;
			{9'd292, 8'd30}: color_data = 12'h660;
			{9'd292, 8'd31}: color_data = 12'h660;
			{9'd292, 8'd32}: color_data = 12'h110;
			{9'd292, 8'd68}: color_data = 12'h047;
			{9'd292, 8'd69}: color_data = 12'h6df;
			{9'd292, 8'd70}: color_data = 12'heff;
			{9'd292, 8'd71}: color_data = 12'h6df;
			{9'd292, 8'd72}: color_data = 12'h0bf;
			{9'd292, 8'd73}: color_data = 12'h0bf;
			{9'd292, 8'd74}: color_data = 12'h056;
			{9'd292, 8'd75}: color_data = 12'h012;
			{9'd292, 8'd76}: color_data = 12'h08b;
			{9'd292, 8'd77}: color_data = 12'h034;
			{9'd292, 8'd128}: color_data = 12'h047;
			{9'd292, 8'd129}: color_data = 12'h6df;
			{9'd292, 8'd130}: color_data = 12'heff;
			{9'd292, 8'd131}: color_data = 12'h6df;
			{9'd292, 8'd132}: color_data = 12'h0bf;
			{9'd292, 8'd133}: color_data = 12'h0bf;
			{9'd292, 8'd134}: color_data = 12'h056;
			{9'd292, 8'd135}: color_data = 12'h012;
			{9'd292, 8'd136}: color_data = 12'h08b;
			{9'd292, 8'd137}: color_data = 12'h034;
			{9'd292, 8'd170}: color_data = 12'h000;
			{9'd292, 8'd171}: color_data = 12'h068;
			{9'd292, 8'd172}: color_data = 12'h8ef;
			{9'd292, 8'd173}: color_data = 12'hdff;
			{9'd292, 8'd174}: color_data = 12'h4cf;
			{9'd292, 8'd175}: color_data = 12'h0cf;
			{9'd292, 8'd176}: color_data = 12'h0ae;
			{9'd292, 8'd177}: color_data = 12'h035;
			{9'd292, 8'd178}: color_data = 12'h023;
			{9'd292, 8'd179}: color_data = 12'h08c;
			{9'd292, 8'd180}: color_data = 12'h023;
			{9'd292, 8'd222}: color_data = 12'h200;
			{9'd292, 8'd223}: color_data = 12'h900;
			{9'd292, 8'd224}: color_data = 12'hb00;
			{9'd292, 8'd225}: color_data = 12'h800;
			{9'd292, 8'd226}: color_data = 12'h200;
			{9'd292, 8'd227}: color_data = 12'hb30;
			{9'd292, 8'd228}: color_data = 12'hc10;
			{9'd292, 8'd229}: color_data = 12'h800;
			{9'd292, 8'd230}: color_data = 12'h300;
			{9'd292, 8'd231}: color_data = 12'h400;
			{9'd292, 8'd232}: color_data = 12'ha00;
			{9'd292, 8'd233}: color_data = 12'ha00;
			{9'd292, 8'd234}: color_data = 12'h500;
			{9'd292, 8'd235}: color_data = 12'h510;
			{9'd292, 8'd236}: color_data = 12'hd30;
			{9'd292, 8'd237}: color_data = 12'ha00;
			{9'd292, 8'd238}: color_data = 12'h700;
			{9'd292, 8'd239}: color_data = 12'h100;
			{9'd293, 8'd16}: color_data = 12'h010;
			{9'd293, 8'd17}: color_data = 12'h780;
			{9'd293, 8'd18}: color_data = 12'hac0;
			{9'd293, 8'd19}: color_data = 12'hdea;
			{9'd293, 8'd20}: color_data = 12'hfff;
			{9'd293, 8'd21}: color_data = 12'hcd7;
			{9'd293, 8'd22}: color_data = 12'h9b0;
			{9'd293, 8'd23}: color_data = 12'h9b0;
			{9'd293, 8'd24}: color_data = 12'h9b0;
			{9'd293, 8'd25}: color_data = 12'h8a0;
			{9'd293, 8'd26}: color_data = 12'h450;
			{9'd293, 8'd27}: color_data = 12'h020;
			{9'd293, 8'd28}: color_data = 12'h140;
			{9'd293, 8'd29}: color_data = 12'h240;
			{9'd293, 8'd30}: color_data = 12'h660;
			{9'd293, 8'd31}: color_data = 12'h660;
			{9'd293, 8'd32}: color_data = 12'h110;
			{9'd293, 8'd68}: color_data = 12'h047;
			{9'd293, 8'd69}: color_data = 12'h6df;
			{9'd293, 8'd70}: color_data = 12'hfff;
			{9'd293, 8'd71}: color_data = 12'hdff;
			{9'd293, 8'd72}: color_data = 12'h5df;
			{9'd293, 8'd73}: color_data = 12'h068;
			{9'd293, 8'd74}: color_data = 12'h000;
			{9'd293, 8'd75}: color_data = 12'h012;
			{9'd293, 8'd76}: color_data = 12'h08c;
			{9'd293, 8'd77}: color_data = 12'h034;
			{9'd293, 8'd128}: color_data = 12'h047;
			{9'd293, 8'd129}: color_data = 12'h6df;
			{9'd293, 8'd130}: color_data = 12'hfff;
			{9'd293, 8'd131}: color_data = 12'hdff;
			{9'd293, 8'd132}: color_data = 12'h5df;
			{9'd293, 8'd133}: color_data = 12'h068;
			{9'd293, 8'd134}: color_data = 12'h000;
			{9'd293, 8'd135}: color_data = 12'h012;
			{9'd293, 8'd136}: color_data = 12'h08c;
			{9'd293, 8'd137}: color_data = 12'h034;
			{9'd293, 8'd170}: color_data = 12'h000;
			{9'd293, 8'd171}: color_data = 12'h068;
			{9'd293, 8'd172}: color_data = 12'h8ef;
			{9'd293, 8'd173}: color_data = 12'hfff;
			{9'd293, 8'd174}: color_data = 12'hcff;
			{9'd293, 8'd175}: color_data = 12'h4ce;
			{9'd293, 8'd176}: color_data = 12'h057;
			{9'd293, 8'd177}: color_data = 12'h000;
			{9'd293, 8'd178}: color_data = 12'h023;
			{9'd293, 8'd179}: color_data = 12'h08c;
			{9'd293, 8'd180}: color_data = 12'h023;
			{9'd293, 8'd222}: color_data = 12'h200;
			{9'd293, 8'd223}: color_data = 12'h900;
			{9'd293, 8'd224}: color_data = 12'ha00;
			{9'd293, 8'd225}: color_data = 12'h700;
			{9'd293, 8'd226}: color_data = 12'h200;
			{9'd293, 8'd227}: color_data = 12'hb30;
			{9'd293, 8'd228}: color_data = 12'he20;
			{9'd293, 8'd229}: color_data = 12'ha00;
			{9'd293, 8'd230}: color_data = 12'h300;
			{9'd293, 8'd231}: color_data = 12'h400;
			{9'd293, 8'd232}: color_data = 12'ha00;
			{9'd293, 8'd233}: color_data = 12'ha00;
			{9'd293, 8'd234}: color_data = 12'h400;
			{9'd293, 8'd235}: color_data = 12'h510;
			{9'd293, 8'd236}: color_data = 12'hf40;
			{9'd293, 8'd237}: color_data = 12'hd10;
			{9'd293, 8'd238}: color_data = 12'h800;
			{9'd293, 8'd239}: color_data = 12'h100;
			{9'd294, 8'd16}: color_data = 12'h010;
			{9'd294, 8'd17}: color_data = 12'h780;
			{9'd294, 8'd18}: color_data = 12'hac0;
			{9'd294, 8'd19}: color_data = 12'hdea;
			{9'd294, 8'd20}: color_data = 12'hfff;
			{9'd294, 8'd21}: color_data = 12'hcd7;
			{9'd294, 8'd22}: color_data = 12'h9b0;
			{9'd294, 8'd23}: color_data = 12'h9b0;
			{9'd294, 8'd24}: color_data = 12'h9b0;
			{9'd294, 8'd25}: color_data = 12'h8a0;
			{9'd294, 8'd26}: color_data = 12'h450;
			{9'd294, 8'd27}: color_data = 12'h020;
			{9'd294, 8'd28}: color_data = 12'h140;
			{9'd294, 8'd29}: color_data = 12'h240;
			{9'd294, 8'd30}: color_data = 12'h660;
			{9'd294, 8'd31}: color_data = 12'h660;
			{9'd294, 8'd32}: color_data = 12'h110;
			{9'd294, 8'd68}: color_data = 12'h047;
			{9'd294, 8'd69}: color_data = 12'h6df;
			{9'd294, 8'd70}: color_data = 12'hfff;
			{9'd294, 8'd71}: color_data = 12'hfff;
			{9'd294, 8'd72}: color_data = 12'h9aa;
			{9'd294, 8'd73}: color_data = 12'h011;
			{9'd294, 8'd75}: color_data = 12'h012;
			{9'd294, 8'd76}: color_data = 12'h08c;
			{9'd294, 8'd77}: color_data = 12'h034;
			{9'd294, 8'd128}: color_data = 12'h047;
			{9'd294, 8'd129}: color_data = 12'h6df;
			{9'd294, 8'd130}: color_data = 12'hfff;
			{9'd294, 8'd131}: color_data = 12'hfff;
			{9'd294, 8'd132}: color_data = 12'h9aa;
			{9'd294, 8'd133}: color_data = 12'h111;
			{9'd294, 8'd135}: color_data = 12'h012;
			{9'd294, 8'd136}: color_data = 12'h08c;
			{9'd294, 8'd137}: color_data = 12'h034;
			{9'd294, 8'd170}: color_data = 12'h000;
			{9'd294, 8'd171}: color_data = 12'h068;
			{9'd294, 8'd172}: color_data = 12'h7ef;
			{9'd294, 8'd173}: color_data = 12'hfff;
			{9'd294, 8'd174}: color_data = 12'hfff;
			{9'd294, 8'd175}: color_data = 12'h899;
			{9'd294, 8'd176}: color_data = 12'h001;
			{9'd294, 8'd178}: color_data = 12'h024;
			{9'd294, 8'd179}: color_data = 12'h08c;
			{9'd294, 8'd180}: color_data = 12'h023;
			{9'd294, 8'd222}: color_data = 12'h200;
			{9'd294, 8'd223}: color_data = 12'h800;
			{9'd294, 8'd224}: color_data = 12'ha00;
			{9'd294, 8'd225}: color_data = 12'h700;
			{9'd294, 8'd226}: color_data = 12'h200;
			{9'd294, 8'd227}: color_data = 12'h920;
			{9'd294, 8'd228}: color_data = 12'hd30;
			{9'd294, 8'd229}: color_data = 12'h910;
			{9'd294, 8'd230}: color_data = 12'h200;
			{9'd294, 8'd231}: color_data = 12'h400;
			{9'd294, 8'd232}: color_data = 12'h900;
			{9'd294, 8'd233}: color_data = 12'ha00;
			{9'd294, 8'd234}: color_data = 12'h400;
			{9'd294, 8'd235}: color_data = 12'h310;
			{9'd294, 8'd236}: color_data = 12'hc30;
			{9'd294, 8'd237}: color_data = 12'hc20;
			{9'd294, 8'd238}: color_data = 12'h600;
			{9'd294, 8'd239}: color_data = 12'h000;
			{9'd295, 8'd16}: color_data = 12'h010;
			{9'd295, 8'd17}: color_data = 12'h780;
			{9'd295, 8'd18}: color_data = 12'hac0;
			{9'd295, 8'd19}: color_data = 12'hdea;
			{9'd295, 8'd20}: color_data = 12'hfff;
			{9'd295, 8'd21}: color_data = 12'hcd7;
			{9'd295, 8'd22}: color_data = 12'h9b0;
			{9'd295, 8'd23}: color_data = 12'h9b0;
			{9'd295, 8'd24}: color_data = 12'h9b0;
			{9'd295, 8'd25}: color_data = 12'h8a0;
			{9'd295, 8'd26}: color_data = 12'h450;
			{9'd295, 8'd27}: color_data = 12'h020;
			{9'd295, 8'd28}: color_data = 12'h140;
			{9'd295, 8'd29}: color_data = 12'h240;
			{9'd295, 8'd30}: color_data = 12'h660;
			{9'd295, 8'd31}: color_data = 12'h660;
			{9'd295, 8'd32}: color_data = 12'h110;
			{9'd295, 8'd68}: color_data = 12'h047;
			{9'd295, 8'd69}: color_data = 12'h6df;
			{9'd295, 8'd70}: color_data = 12'hfff;
			{9'd295, 8'd71}: color_data = 12'hcbb;
			{9'd295, 8'd72}: color_data = 12'h323;
			{9'd295, 8'd73}: color_data = 12'h002;
			{9'd295, 8'd74}: color_data = 12'h000;
			{9'd295, 8'd75}: color_data = 12'h012;
			{9'd295, 8'd76}: color_data = 12'h08c;
			{9'd295, 8'd77}: color_data = 12'h034;
			{9'd295, 8'd128}: color_data = 12'h047;
			{9'd295, 8'd129}: color_data = 12'h6df;
			{9'd295, 8'd130}: color_data = 12'hfff;
			{9'd295, 8'd131}: color_data = 12'hcbb;
			{9'd295, 8'd132}: color_data = 12'h323;
			{9'd295, 8'd133}: color_data = 12'h002;
			{9'd295, 8'd134}: color_data = 12'h000;
			{9'd295, 8'd135}: color_data = 12'h012;
			{9'd295, 8'd136}: color_data = 12'h08c;
			{9'd295, 8'd137}: color_data = 12'h034;
			{9'd295, 8'd170}: color_data = 12'h000;
			{9'd295, 8'd171}: color_data = 12'h068;
			{9'd295, 8'd172}: color_data = 12'h8ef;
			{9'd295, 8'd173}: color_data = 12'hfff;
			{9'd295, 8'd174}: color_data = 12'haaa;
			{9'd295, 8'd175}: color_data = 12'h212;
			{9'd295, 8'd176}: color_data = 12'h002;
			{9'd295, 8'd178}: color_data = 12'h023;
			{9'd295, 8'd179}: color_data = 12'h08c;
			{9'd295, 8'd180}: color_data = 12'h023;
			{9'd295, 8'd222}: color_data = 12'h200;
			{9'd295, 8'd223}: color_data = 12'h900;
			{9'd295, 8'd224}: color_data = 12'ha00;
			{9'd295, 8'd225}: color_data = 12'h800;
			{9'd295, 8'd226}: color_data = 12'h100;
			{9'd295, 8'd227}: color_data = 12'h100;
			{9'd295, 8'd228}: color_data = 12'h310;
			{9'd295, 8'd229}: color_data = 12'h200;
			{9'd295, 8'd230}: color_data = 12'h000;
			{9'd295, 8'd231}: color_data = 12'h500;
			{9'd295, 8'd232}: color_data = 12'ha00;
			{9'd295, 8'd233}: color_data = 12'ha00;
			{9'd295, 8'd234}: color_data = 12'h500;
			{9'd295, 8'd235}: color_data = 12'h000;
			{9'd295, 8'd236}: color_data = 12'h200;
			{9'd295, 8'd237}: color_data = 12'h300;
			{9'd295, 8'd238}: color_data = 12'h100;
			{9'd295, 8'd239}: color_data = 12'h000;
			{9'd296, 8'd16}: color_data = 12'h010;
			{9'd296, 8'd17}: color_data = 12'h780;
			{9'd296, 8'd18}: color_data = 12'hac0;
			{9'd296, 8'd19}: color_data = 12'hdea;
			{9'd296, 8'd20}: color_data = 12'hfff;
			{9'd296, 8'd21}: color_data = 12'hcd7;
			{9'd296, 8'd22}: color_data = 12'h9b0;
			{9'd296, 8'd23}: color_data = 12'h9b0;
			{9'd296, 8'd24}: color_data = 12'h9b0;
			{9'd296, 8'd25}: color_data = 12'h8a0;
			{9'd296, 8'd26}: color_data = 12'h450;
			{9'd296, 8'd27}: color_data = 12'h020;
			{9'd296, 8'd28}: color_data = 12'h140;
			{9'd296, 8'd29}: color_data = 12'h240;
			{9'd296, 8'd30}: color_data = 12'h660;
			{9'd296, 8'd31}: color_data = 12'h660;
			{9'd296, 8'd32}: color_data = 12'h110;
			{9'd296, 8'd68}: color_data = 12'h047;
			{9'd296, 8'd69}: color_data = 12'h6ef;
			{9'd296, 8'd70}: color_data = 12'hdcc;
			{9'd296, 8'd71}: color_data = 12'h434;
			{9'd296, 8'd72}: color_data = 12'h003;
			{9'd296, 8'd73}: color_data = 12'h005;
			{9'd296, 8'd74}: color_data = 12'h002;
			{9'd296, 8'd75}: color_data = 12'h012;
			{9'd296, 8'd76}: color_data = 12'h08c;
			{9'd296, 8'd77}: color_data = 12'h034;
			{9'd296, 8'd128}: color_data = 12'h047;
			{9'd296, 8'd129}: color_data = 12'h6ef;
			{9'd296, 8'd130}: color_data = 12'hddc;
			{9'd296, 8'd131}: color_data = 12'h434;
			{9'd296, 8'd132}: color_data = 12'h003;
			{9'd296, 8'd133}: color_data = 12'h005;
			{9'd296, 8'd134}: color_data = 12'h002;
			{9'd296, 8'd135}: color_data = 12'h012;
			{9'd296, 8'd136}: color_data = 12'h08c;
			{9'd296, 8'd137}: color_data = 12'h034;
			{9'd296, 8'd170}: color_data = 12'h000;
			{9'd296, 8'd171}: color_data = 12'h068;
			{9'd296, 8'd172}: color_data = 12'h8ff;
			{9'd296, 8'd173}: color_data = 12'hcbb;
			{9'd296, 8'd174}: color_data = 12'h323;
			{9'd296, 8'd175}: color_data = 12'h003;
			{9'd296, 8'd176}: color_data = 12'h005;
			{9'd296, 8'd177}: color_data = 12'h002;
			{9'd296, 8'd178}: color_data = 12'h023;
			{9'd296, 8'd179}: color_data = 12'h09c;
			{9'd296, 8'd180}: color_data = 12'h023;
			{9'd296, 8'd222}: color_data = 12'h300;
			{9'd296, 8'd223}: color_data = 12'hc20;
			{9'd296, 8'd224}: color_data = 12'ha00;
			{9'd296, 8'd225}: color_data = 12'h800;
			{9'd296, 8'd226}: color_data = 12'h100;
			{9'd296, 8'd227}: color_data = 12'h300;
			{9'd296, 8'd228}: color_data = 12'h500;
			{9'd296, 8'd229}: color_data = 12'h500;
			{9'd296, 8'd230}: color_data = 12'h100;
			{9'd296, 8'd231}: color_data = 12'h710;
			{9'd296, 8'd232}: color_data = 12'hc10;
			{9'd296, 8'd233}: color_data = 12'h900;
			{9'd296, 8'd234}: color_data = 12'h500;
			{9'd296, 8'd235}: color_data = 12'h100;
			{9'd296, 8'd236}: color_data = 12'h500;
			{9'd296, 8'd237}: color_data = 12'h600;
			{9'd296, 8'd238}: color_data = 12'h400;
			{9'd296, 8'd239}: color_data = 12'h000;
			{9'd297, 8'd16}: color_data = 12'h010;
			{9'd297, 8'd17}: color_data = 12'h780;
			{9'd297, 8'd18}: color_data = 12'hac0;
			{9'd297, 8'd19}: color_data = 12'hdea;
			{9'd297, 8'd20}: color_data = 12'hfff;
			{9'd297, 8'd21}: color_data = 12'hcd7;
			{9'd297, 8'd22}: color_data = 12'h9b0;
			{9'd297, 8'd23}: color_data = 12'h9b0;
			{9'd297, 8'd24}: color_data = 12'h9b0;
			{9'd297, 8'd25}: color_data = 12'h8a0;
			{9'd297, 8'd26}: color_data = 12'h450;
			{9'd297, 8'd27}: color_data = 12'h020;
			{9'd297, 8'd28}: color_data = 12'h140;
			{9'd297, 8'd29}: color_data = 12'h240;
			{9'd297, 8'd30}: color_data = 12'h660;
			{9'd297, 8'd31}: color_data = 12'h660;
			{9'd297, 8'd32}: color_data = 12'h110;
			{9'd297, 8'd68}: color_data = 12'h057;
			{9'd297, 8'd69}: color_data = 12'h3bd;
			{9'd297, 8'd70}: color_data = 12'h555;
			{9'd297, 8'd71}: color_data = 12'h002;
			{9'd297, 8'd72}: color_data = 12'h005;
			{9'd297, 8'd73}: color_data = 12'h005;
			{9'd297, 8'd74}: color_data = 12'h004;
			{9'd297, 8'd75}: color_data = 12'h025;
			{9'd297, 8'd76}: color_data = 12'h09c;
			{9'd297, 8'd77}: color_data = 12'h034;
			{9'd297, 8'd128}: color_data = 12'h057;
			{9'd297, 8'd129}: color_data = 12'h3bd;
			{9'd297, 8'd130}: color_data = 12'h555;
			{9'd297, 8'd131}: color_data = 12'h002;
			{9'd297, 8'd132}: color_data = 12'h005;
			{9'd297, 8'd133}: color_data = 12'h005;
			{9'd297, 8'd134}: color_data = 12'h004;
			{9'd297, 8'd135}: color_data = 12'h025;
			{9'd297, 8'd136}: color_data = 12'h09c;
			{9'd297, 8'd137}: color_data = 12'h034;
			{9'd297, 8'd170}: color_data = 12'h000;
			{9'd297, 8'd171}: color_data = 12'h079;
			{9'd297, 8'd172}: color_data = 12'h4bd;
			{9'd297, 8'd173}: color_data = 12'h444;
			{9'd297, 8'd174}: color_data = 12'h002;
			{9'd297, 8'd175}: color_data = 12'h005;
			{9'd297, 8'd176}: color_data = 12'h005;
			{9'd297, 8'd177}: color_data = 12'h004;
			{9'd297, 8'd178}: color_data = 12'h036;
			{9'd297, 8'd179}: color_data = 12'h09c;
			{9'd297, 8'd180}: color_data = 12'h023;
			{9'd297, 8'd222}: color_data = 12'h410;
			{9'd297, 8'd223}: color_data = 12'hd30;
			{9'd297, 8'd224}: color_data = 12'hb00;
			{9'd297, 8'd225}: color_data = 12'h700;
			{9'd297, 8'd226}: color_data = 12'h200;
			{9'd297, 8'd227}: color_data = 12'h700;
			{9'd297, 8'd228}: color_data = 12'hb00;
			{9'd297, 8'd229}: color_data = 12'h900;
			{9'd297, 8'd230}: color_data = 12'h300;
			{9'd297, 8'd231}: color_data = 12'h820;
			{9'd297, 8'd232}: color_data = 12'hd20;
			{9'd297, 8'd233}: color_data = 12'h900;
			{9'd297, 8'd234}: color_data = 12'h500;
			{9'd297, 8'd235}: color_data = 12'h300;
			{9'd297, 8'd236}: color_data = 12'h900;
			{9'd297, 8'd237}: color_data = 12'hb00;
			{9'd297, 8'd238}: color_data = 12'h800;
			{9'd297, 8'd239}: color_data = 12'h100;
			{9'd298, 8'd16}: color_data = 12'h010;
			{9'd298, 8'd17}: color_data = 12'h780;
			{9'd298, 8'd18}: color_data = 12'hac0;
			{9'd298, 8'd19}: color_data = 12'hdea;
			{9'd298, 8'd20}: color_data = 12'hfff;
			{9'd298, 8'd21}: color_data = 12'hcd7;
			{9'd298, 8'd22}: color_data = 12'h9b0;
			{9'd298, 8'd23}: color_data = 12'h9b0;
			{9'd298, 8'd24}: color_data = 12'h9b0;
			{9'd298, 8'd25}: color_data = 12'h8a0;
			{9'd298, 8'd26}: color_data = 12'h450;
			{9'd298, 8'd27}: color_data = 12'h020;
			{9'd298, 8'd28}: color_data = 12'h140;
			{9'd298, 8'd29}: color_data = 12'h240;
			{9'd298, 8'd30}: color_data = 12'h660;
			{9'd298, 8'd31}: color_data = 12'h660;
			{9'd298, 8'd32}: color_data = 12'h110;
			{9'd298, 8'd68}: color_data = 12'h035;
			{9'd298, 8'd69}: color_data = 12'h047;
			{9'd298, 8'd70}: color_data = 12'h001;
			{9'd298, 8'd71}: color_data = 12'h004;
			{9'd298, 8'd72}: color_data = 12'h004;
			{9'd298, 8'd73}: color_data = 12'h004;
			{9'd298, 8'd74}: color_data = 12'h004;
			{9'd298, 8'd75}: color_data = 12'h015;
			{9'd298, 8'd76}: color_data = 12'h059;
			{9'd298, 8'd77}: color_data = 12'h023;
			{9'd298, 8'd128}: color_data = 12'h035;
			{9'd298, 8'd129}: color_data = 12'h047;
			{9'd298, 8'd130}: color_data = 12'h001;
			{9'd298, 8'd131}: color_data = 12'h004;
			{9'd298, 8'd132}: color_data = 12'h004;
			{9'd298, 8'd133}: color_data = 12'h004;
			{9'd298, 8'd134}: color_data = 12'h004;
			{9'd298, 8'd135}: color_data = 12'h015;
			{9'd298, 8'd136}: color_data = 12'h059;
			{9'd298, 8'd137}: color_data = 12'h023;
			{9'd298, 8'd170}: color_data = 12'h000;
			{9'd298, 8'd171}: color_data = 12'h047;
			{9'd298, 8'd172}: color_data = 12'h036;
			{9'd298, 8'd173}: color_data = 12'h001;
			{9'd298, 8'd174}: color_data = 12'h004;
			{9'd298, 8'd175}: color_data = 12'h004;
			{9'd298, 8'd176}: color_data = 12'h004;
			{9'd298, 8'd177}: color_data = 12'h004;
			{9'd298, 8'd178}: color_data = 12'h016;
			{9'd298, 8'd179}: color_data = 12'h059;
			{9'd298, 8'd180}: color_data = 12'h012;
			{9'd298, 8'd222}: color_data = 12'h410;
			{9'd298, 8'd223}: color_data = 12'he40;
			{9'd298, 8'd224}: color_data = 12'hd20;
			{9'd298, 8'd225}: color_data = 12'h800;
			{9'd298, 8'd226}: color_data = 12'h200;
			{9'd298, 8'd227}: color_data = 12'h600;
			{9'd298, 8'd228}: color_data = 12'ha00;
			{9'd298, 8'd229}: color_data = 12'h900;
			{9'd298, 8'd230}: color_data = 12'h300;
			{9'd298, 8'd231}: color_data = 12'h820;
			{9'd298, 8'd232}: color_data = 12'hf30;
			{9'd298, 8'd233}: color_data = 12'hc00;
			{9'd298, 8'd234}: color_data = 12'h500;
			{9'd298, 8'd235}: color_data = 12'h200;
			{9'd298, 8'd236}: color_data = 12'h900;
			{9'd298, 8'd237}: color_data = 12'ha00;
			{9'd298, 8'd238}: color_data = 12'h700;
			{9'd298, 8'd239}: color_data = 12'h100;
			{9'd299, 8'd16}: color_data = 12'h010;
			{9'd299, 8'd17}: color_data = 12'h780;
			{9'd299, 8'd18}: color_data = 12'hac0;
			{9'd299, 8'd19}: color_data = 12'hdea;
			{9'd299, 8'd20}: color_data = 12'hfff;
			{9'd299, 8'd21}: color_data = 12'hcd7;
			{9'd299, 8'd22}: color_data = 12'h9b0;
			{9'd299, 8'd23}: color_data = 12'h9b0;
			{9'd299, 8'd24}: color_data = 12'h9b0;
			{9'd299, 8'd25}: color_data = 12'h8a0;
			{9'd299, 8'd26}: color_data = 12'h450;
			{9'd299, 8'd27}: color_data = 12'h020;
			{9'd299, 8'd28}: color_data = 12'h140;
			{9'd299, 8'd29}: color_data = 12'h240;
			{9'd299, 8'd30}: color_data = 12'h660;
			{9'd299, 8'd31}: color_data = 12'h660;
			{9'd299, 8'd32}: color_data = 12'h220;
			{9'd299, 8'd33}: color_data = 12'h000;
			{9'd299, 8'd45}: color_data = 12'h000;
			{9'd299, 8'd46}: color_data = 12'h110;
			{9'd299, 8'd47}: color_data = 12'h110;
			{9'd299, 8'd48}: color_data = 12'h110;
			{9'd299, 8'd49}: color_data = 12'h110;
			{9'd299, 8'd50}: color_data = 12'h000;
			{9'd299, 8'd68}: color_data = 12'h013;
			{9'd299, 8'd69}: color_data = 12'h027;
			{9'd299, 8'd70}: color_data = 12'h016;
			{9'd299, 8'd71}: color_data = 12'h027;
			{9'd299, 8'd72}: color_data = 12'h027;
			{9'd299, 8'd73}: color_data = 12'h027;
			{9'd299, 8'd74}: color_data = 12'h027;
			{9'd299, 8'd75}: color_data = 12'h028;
			{9'd299, 8'd76}: color_data = 12'h027;
			{9'd299, 8'd77}: color_data = 12'h001;
			{9'd299, 8'd128}: color_data = 12'h013;
			{9'd299, 8'd129}: color_data = 12'h027;
			{9'd299, 8'd130}: color_data = 12'h016;
			{9'd299, 8'd131}: color_data = 12'h027;
			{9'd299, 8'd132}: color_data = 12'h027;
			{9'd299, 8'd133}: color_data = 12'h027;
			{9'd299, 8'd134}: color_data = 12'h027;
			{9'd299, 8'd135}: color_data = 12'h028;
			{9'd299, 8'd136}: color_data = 12'h027;
			{9'd299, 8'd137}: color_data = 12'h001;
			{9'd299, 8'd170}: color_data = 12'h000;
			{9'd299, 8'd171}: color_data = 12'h014;
			{9'd299, 8'd172}: color_data = 12'h027;
			{9'd299, 8'd173}: color_data = 12'h016;
			{9'd299, 8'd174}: color_data = 12'h027;
			{9'd299, 8'd175}: color_data = 12'h027;
			{9'd299, 8'd176}: color_data = 12'h027;
			{9'd299, 8'd177}: color_data = 12'h027;
			{9'd299, 8'd178}: color_data = 12'h028;
			{9'd299, 8'd179}: color_data = 12'h026;
			{9'd299, 8'd180}: color_data = 12'h001;
			{9'd299, 8'd204}: color_data = 12'h000;
			{9'd299, 8'd205}: color_data = 12'h221;
			{9'd299, 8'd206}: color_data = 12'h333;
			{9'd299, 8'd207}: color_data = 12'h222;
			{9'd299, 8'd208}: color_data = 12'h333;
			{9'd299, 8'd209}: color_data = 12'h323;
			{9'd299, 8'd210}: color_data = 12'h120;
			{9'd299, 8'd211}: color_data = 12'h120;
			{9'd299, 8'd212}: color_data = 12'h120;
			{9'd299, 8'd213}: color_data = 12'h120;
			{9'd299, 8'd214}: color_data = 12'h120;
			{9'd299, 8'd215}: color_data = 12'h110;
			{9'd299, 8'd216}: color_data = 12'h000;
			{9'd299, 8'd217}: color_data = 12'h000;
			{9'd299, 8'd218}: color_data = 12'h000;
			{9'd299, 8'd219}: color_data = 12'h000;
			{9'd299, 8'd220}: color_data = 12'h110;
			{9'd299, 8'd221}: color_data = 12'h000;
			{9'd299, 8'd222}: color_data = 12'h200;
			{9'd299, 8'd223}: color_data = 12'hb30;
			{9'd299, 8'd224}: color_data = 12'hc30;
			{9'd299, 8'd225}: color_data = 12'h700;
			{9'd299, 8'd226}: color_data = 12'h100;
			{9'd299, 8'd227}: color_data = 12'h600;
			{9'd299, 8'd228}: color_data = 12'ha00;
			{9'd299, 8'd229}: color_data = 12'h900;
			{9'd299, 8'd230}: color_data = 12'h300;
			{9'd299, 8'd231}: color_data = 12'h620;
			{9'd299, 8'd232}: color_data = 12'hd40;
			{9'd299, 8'd233}: color_data = 12'ha20;
			{9'd299, 8'd234}: color_data = 12'h300;
			{9'd299, 8'd235}: color_data = 12'h200;
			{9'd299, 8'd236}: color_data = 12'h800;
			{9'd299, 8'd237}: color_data = 12'ha00;
			{9'd299, 8'd238}: color_data = 12'h700;
			{9'd299, 8'd239}: color_data = 12'h100;
			{9'd300, 8'd16}: color_data = 12'h010;
			{9'd300, 8'd17}: color_data = 12'h780;
			{9'd300, 8'd18}: color_data = 12'hac0;
			{9'd300, 8'd19}: color_data = 12'hdea;
			{9'd300, 8'd20}: color_data = 12'hfff;
			{9'd300, 8'd21}: color_data = 12'hcd7;
			{9'd300, 8'd22}: color_data = 12'h9b0;
			{9'd300, 8'd23}: color_data = 12'h9b0;
			{9'd300, 8'd24}: color_data = 12'h9b0;
			{9'd300, 8'd25}: color_data = 12'h8a0;
			{9'd300, 8'd26}: color_data = 12'h450;
			{9'd300, 8'd27}: color_data = 12'h020;
			{9'd300, 8'd28}: color_data = 12'h140;
			{9'd300, 8'd29}: color_data = 12'h240;
			{9'd300, 8'd30}: color_data = 12'h560;
			{9'd300, 8'd31}: color_data = 12'h660;
			{9'd300, 8'd32}: color_data = 12'h550;
			{9'd300, 8'd33}: color_data = 12'h110;
			{9'd300, 8'd34}: color_data = 12'h000;
			{9'd300, 8'd35}: color_data = 12'h000;
			{9'd300, 8'd36}: color_data = 12'h000;
			{9'd300, 8'd37}: color_data = 12'h000;
			{9'd300, 8'd38}: color_data = 12'h000;
			{9'd300, 8'd39}: color_data = 12'h000;
			{9'd300, 8'd40}: color_data = 12'h000;
			{9'd300, 8'd41}: color_data = 12'h000;
			{9'd300, 8'd42}: color_data = 12'h000;
			{9'd300, 8'd43}: color_data = 12'h000;
			{9'd300, 8'd44}: color_data = 12'h000;
			{9'd300, 8'd45}: color_data = 12'h110;
			{9'd300, 8'd46}: color_data = 12'h670;
			{9'd300, 8'd47}: color_data = 12'h670;
			{9'd300, 8'd48}: color_data = 12'h550;
			{9'd300, 8'd49}: color_data = 12'h550;
			{9'd300, 8'd50}: color_data = 12'h220;
			{9'd300, 8'd51}: color_data = 12'h000;
			{9'd300, 8'd52}: color_data = 12'h000;
			{9'd300, 8'd53}: color_data = 12'h000;
			{9'd300, 8'd54}: color_data = 12'h000;
			{9'd300, 8'd55}: color_data = 12'h000;
			{9'd300, 8'd56}: color_data = 12'h000;
			{9'd300, 8'd57}: color_data = 12'h000;
			{9'd300, 8'd68}: color_data = 12'h035;
			{9'd300, 8'd69}: color_data = 12'h09e;
			{9'd300, 8'd70}: color_data = 12'h09e;
			{9'd300, 8'd71}: color_data = 12'h09e;
			{9'd300, 8'd72}: color_data = 12'h09e;
			{9'd300, 8'd73}: color_data = 12'h09e;
			{9'd300, 8'd74}: color_data = 12'h09e;
			{9'd300, 8'd75}: color_data = 12'h09e;
			{9'd300, 8'd76}: color_data = 12'h08c;
			{9'd300, 8'd77}: color_data = 12'h023;
			{9'd300, 8'd128}: color_data = 12'h035;
			{9'd300, 8'd129}: color_data = 12'h09e;
			{9'd300, 8'd130}: color_data = 12'h09e;
			{9'd300, 8'd131}: color_data = 12'h09e;
			{9'd300, 8'd132}: color_data = 12'h09e;
			{9'd300, 8'd133}: color_data = 12'h09e;
			{9'd300, 8'd134}: color_data = 12'h09e;
			{9'd300, 8'd135}: color_data = 12'h09e;
			{9'd300, 8'd136}: color_data = 12'h08c;
			{9'd300, 8'd137}: color_data = 12'h023;
			{9'd300, 8'd170}: color_data = 12'h000;
			{9'd300, 8'd171}: color_data = 12'h057;
			{9'd300, 8'd172}: color_data = 12'h0ae;
			{9'd300, 8'd173}: color_data = 12'h09e;
			{9'd300, 8'd174}: color_data = 12'h09e;
			{9'd300, 8'd175}: color_data = 12'h09e;
			{9'd300, 8'd176}: color_data = 12'h09e;
			{9'd300, 8'd177}: color_data = 12'h09e;
			{9'd300, 8'd178}: color_data = 12'h09e;
			{9'd300, 8'd179}: color_data = 12'h07b;
			{9'd300, 8'd180}: color_data = 12'h012;
			{9'd300, 8'd204}: color_data = 12'h230;
			{9'd300, 8'd205}: color_data = 12'h9b4;
			{9'd300, 8'd206}: color_data = 12'hddc;
			{9'd300, 8'd207}: color_data = 12'hddd;
			{9'd300, 8'd208}: color_data = 12'hddd;
			{9'd300, 8'd209}: color_data = 12'hccb;
			{9'd300, 8'd210}: color_data = 12'h8a1;
			{9'd300, 8'd211}: color_data = 12'h790;
			{9'd300, 8'd212}: color_data = 12'h790;
			{9'd300, 8'd213}: color_data = 12'h890;
			{9'd300, 8'd214}: color_data = 12'h890;
			{9'd300, 8'd215}: color_data = 12'h670;
			{9'd300, 8'd216}: color_data = 12'h230;
			{9'd300, 8'd217}: color_data = 12'h020;
			{9'd300, 8'd218}: color_data = 12'h130;
			{9'd300, 8'd219}: color_data = 12'h340;
			{9'd300, 8'd220}: color_data = 12'h550;
			{9'd300, 8'd221}: color_data = 12'h330;
			{9'd300, 8'd222}: color_data = 12'h000;
			{9'd300, 8'd223}: color_data = 12'h200;
			{9'd300, 8'd224}: color_data = 12'h300;
			{9'd300, 8'd225}: color_data = 12'h100;
			{9'd300, 8'd226}: color_data = 12'h000;
			{9'd300, 8'd227}: color_data = 12'h700;
			{9'd300, 8'd228}: color_data = 12'ha00;
			{9'd300, 8'd229}: color_data = 12'h900;
			{9'd300, 8'd230}: color_data = 12'h300;
			{9'd300, 8'd231}: color_data = 12'h100;
			{9'd300, 8'd232}: color_data = 12'h310;
			{9'd300, 8'd233}: color_data = 12'h200;
			{9'd300, 8'd234}: color_data = 12'h000;
			{9'd300, 8'd235}: color_data = 12'h300;
			{9'd300, 8'd236}: color_data = 12'h900;
			{9'd300, 8'd237}: color_data = 12'ha00;
			{9'd300, 8'd238}: color_data = 12'h700;
			{9'd300, 8'd239}: color_data = 12'h100;
			{9'd301, 8'd16}: color_data = 12'h010;
			{9'd301, 8'd17}: color_data = 12'h780;
			{9'd301, 8'd18}: color_data = 12'hac0;
			{9'd301, 8'd19}: color_data = 12'hdea;
			{9'd301, 8'd20}: color_data = 12'hfff;
			{9'd301, 8'd21}: color_data = 12'hcd7;
			{9'd301, 8'd22}: color_data = 12'h9b0;
			{9'd301, 8'd23}: color_data = 12'h9b0;
			{9'd301, 8'd24}: color_data = 12'h9b0;
			{9'd301, 8'd25}: color_data = 12'h8a0;
			{9'd301, 8'd26}: color_data = 12'h450;
			{9'd301, 8'd27}: color_data = 12'h020;
			{9'd301, 8'd28}: color_data = 12'h140;
			{9'd301, 8'd29}: color_data = 12'h240;
			{9'd301, 8'd30}: color_data = 12'h350;
			{9'd301, 8'd31}: color_data = 12'h660;
			{9'd301, 8'd32}: color_data = 12'h760;
			{9'd301, 8'd33}: color_data = 12'h550;
			{9'd301, 8'd34}: color_data = 12'h440;
			{9'd301, 8'd35}: color_data = 12'h440;
			{9'd301, 8'd36}: color_data = 12'h440;
			{9'd301, 8'd37}: color_data = 12'h440;
			{9'd301, 8'd38}: color_data = 12'h440;
			{9'd301, 8'd39}: color_data = 12'h440;
			{9'd301, 8'd40}: color_data = 12'h440;
			{9'd301, 8'd41}: color_data = 12'h440;
			{9'd301, 8'd42}: color_data = 12'h440;
			{9'd301, 8'd43}: color_data = 12'h440;
			{9'd301, 8'd44}: color_data = 12'h440;
			{9'd301, 8'd45}: color_data = 12'h550;
			{9'd301, 8'd46}: color_data = 12'h8a0;
			{9'd301, 8'd47}: color_data = 12'h880;
			{9'd301, 8'd48}: color_data = 12'h760;
			{9'd301, 8'd49}: color_data = 12'h770;
			{9'd301, 8'd50}: color_data = 12'h230;
			{9'd301, 8'd51}: color_data = 12'h220;
			{9'd301, 8'd52}: color_data = 12'h440;
			{9'd301, 8'd53}: color_data = 12'h440;
			{9'd301, 8'd54}: color_data = 12'h440;
			{9'd301, 8'd55}: color_data = 12'h440;
			{9'd301, 8'd56}: color_data = 12'h440;
			{9'd301, 8'd57}: color_data = 12'h330;
			{9'd301, 8'd58}: color_data = 12'h000;
			{9'd301, 8'd60}: color_data = 12'h000;
			{9'd301, 8'd68}: color_data = 12'h057;
			{9'd301, 8'd69}: color_data = 12'h4ef;
			{9'd301, 8'd70}: color_data = 12'h7ef;
			{9'd301, 8'd71}: color_data = 12'h0cf;
			{9'd301, 8'd72}: color_data = 12'h0cf;
			{9'd301, 8'd73}: color_data = 12'h0df;
			{9'd301, 8'd74}: color_data = 12'h0bd;
			{9'd301, 8'd75}: color_data = 12'h068;
			{9'd301, 8'd76}: color_data = 12'h09c;
			{9'd301, 8'd77}: color_data = 12'h034;
			{9'd301, 8'd128}: color_data = 12'h057;
			{9'd301, 8'd129}: color_data = 12'h4ef;
			{9'd301, 8'd130}: color_data = 12'h7ef;
			{9'd301, 8'd131}: color_data = 12'h0cf;
			{9'd301, 8'd132}: color_data = 12'h0cf;
			{9'd301, 8'd133}: color_data = 12'h0df;
			{9'd301, 8'd134}: color_data = 12'h0bd;
			{9'd301, 8'd135}: color_data = 12'h068;
			{9'd301, 8'd136}: color_data = 12'h09c;
			{9'd301, 8'd137}: color_data = 12'h034;
			{9'd301, 8'd170}: color_data = 12'h000;
			{9'd301, 8'd171}: color_data = 12'h069;
			{9'd301, 8'd172}: color_data = 12'h6ef;
			{9'd301, 8'd173}: color_data = 12'h6ef;
			{9'd301, 8'd174}: color_data = 12'h0cf;
			{9'd301, 8'd175}: color_data = 12'h0cf;
			{9'd301, 8'd176}: color_data = 12'h0df;
			{9'd301, 8'd177}: color_data = 12'h0ac;
			{9'd301, 8'd178}: color_data = 12'h079;
			{9'd301, 8'd179}: color_data = 12'h09c;
			{9'd301, 8'd180}: color_data = 12'h023;
			{9'd301, 8'd204}: color_data = 12'h340;
			{9'd301, 8'd205}: color_data = 12'had1;
			{9'd301, 8'd206}: color_data = 12'hde9;
			{9'd301, 8'd207}: color_data = 12'hfff;
			{9'd301, 8'd208}: color_data = 12'hffe;
			{9'd301, 8'd209}: color_data = 12'hce6;
			{9'd301, 8'd210}: color_data = 12'hac0;
			{9'd301, 8'd211}: color_data = 12'h9c0;
			{9'd301, 8'd212}: color_data = 12'hac0;
			{9'd301, 8'd213}: color_data = 12'hac0;
			{9'd301, 8'd214}: color_data = 12'hac0;
			{9'd301, 8'd215}: color_data = 12'h890;
			{9'd301, 8'd216}: color_data = 12'h230;
			{9'd301, 8'd217}: color_data = 12'h030;
			{9'd301, 8'd218}: color_data = 12'h140;
			{9'd301, 8'd219}: color_data = 12'h450;
			{9'd301, 8'd220}: color_data = 12'h770;
			{9'd301, 8'd221}: color_data = 12'h450;
			{9'd301, 8'd222}: color_data = 12'h100;
			{9'd301, 8'd223}: color_data = 12'h400;
			{9'd301, 8'd224}: color_data = 12'h600;
			{9'd301, 8'd225}: color_data = 12'h400;
			{9'd301, 8'd226}: color_data = 12'h200;
			{9'd301, 8'd227}: color_data = 12'ha20;
			{9'd301, 8'd228}: color_data = 12'hb10;
			{9'd301, 8'd229}: color_data = 12'h900;
			{9'd301, 8'd230}: color_data = 12'h300;
			{9'd301, 8'd231}: color_data = 12'h200;
			{9'd301, 8'd232}: color_data = 12'h500;
			{9'd301, 8'd233}: color_data = 12'h500;
			{9'd301, 8'd234}: color_data = 12'h200;
			{9'd301, 8'd235}: color_data = 12'h410;
			{9'd301, 8'd236}: color_data = 12'hc20;
			{9'd301, 8'd237}: color_data = 12'ha00;
			{9'd301, 8'd238}: color_data = 12'h700;
			{9'd301, 8'd239}: color_data = 12'h100;
			{9'd302, 8'd16}: color_data = 12'h010;
			{9'd302, 8'd17}: color_data = 12'h780;
			{9'd302, 8'd18}: color_data = 12'hac0;
			{9'd302, 8'd19}: color_data = 12'hdea;
			{9'd302, 8'd20}: color_data = 12'hfff;
			{9'd302, 8'd21}: color_data = 12'hcd7;
			{9'd302, 8'd22}: color_data = 12'h9b0;
			{9'd302, 8'd23}: color_data = 12'h9b0;
			{9'd302, 8'd24}: color_data = 12'h9b0;
			{9'd302, 8'd25}: color_data = 12'h8a0;
			{9'd302, 8'd26}: color_data = 12'h440;
			{9'd302, 8'd27}: color_data = 12'h020;
			{9'd302, 8'd28}: color_data = 12'h140;
			{9'd302, 8'd29}: color_data = 12'h240;
			{9'd302, 8'd30}: color_data = 12'h140;
			{9'd302, 8'd31}: color_data = 12'h350;
			{9'd302, 8'd32}: color_data = 12'h660;
			{9'd302, 8'd33}: color_data = 12'h770;
			{9'd302, 8'd34}: color_data = 12'h670;
			{9'd302, 8'd35}: color_data = 12'h950;
			{9'd302, 8'd36}: color_data = 12'hc30;
			{9'd302, 8'd37}: color_data = 12'hc30;
			{9'd302, 8'd38}: color_data = 12'hc30;
			{9'd302, 8'd39}: color_data = 12'hc30;
			{9'd302, 8'd40}: color_data = 12'hc30;
			{9'd302, 8'd41}: color_data = 12'hc30;
			{9'd302, 8'd42}: color_data = 12'ha40;
			{9'd302, 8'd43}: color_data = 12'h670;
			{9'd302, 8'd44}: color_data = 12'h670;
			{9'd302, 8'd45}: color_data = 12'h770;
			{9'd302, 8'd46}: color_data = 12'h8a0;
			{9'd302, 8'd47}: color_data = 12'h570;
			{9'd302, 8'd48}: color_data = 12'h450;
			{9'd302, 8'd49}: color_data = 12'h450;
			{9'd302, 8'd50}: color_data = 12'h130;
			{9'd302, 8'd51}: color_data = 12'h340;
			{9'd302, 8'd52}: color_data = 12'h770;
			{9'd302, 8'd53}: color_data = 12'h770;
			{9'd302, 8'd54}: color_data = 12'h770;
			{9'd302, 8'd55}: color_data = 12'h770;
			{9'd302, 8'd56}: color_data = 12'h770;
			{9'd302, 8'd57}: color_data = 12'h660;
			{9'd302, 8'd58}: color_data = 12'h330;
			{9'd302, 8'd59}: color_data = 12'h330;
			{9'd302, 8'd60}: color_data = 12'h220;
			{9'd302, 8'd61}: color_data = 12'h000;
			{9'd302, 8'd68}: color_data = 12'h047;
			{9'd302, 8'd69}: color_data = 12'h6df;
			{9'd302, 8'd70}: color_data = 12'heff;
			{9'd302, 8'd71}: color_data = 12'h6df;
			{9'd302, 8'd72}: color_data = 12'h0bf;
			{9'd302, 8'd73}: color_data = 12'h0be;
			{9'd302, 8'd74}: color_data = 12'h056;
			{9'd302, 8'd75}: color_data = 12'h012;
			{9'd302, 8'd76}: color_data = 12'h08b;
			{9'd302, 8'd77}: color_data = 12'h034;
			{9'd302, 8'd128}: color_data = 12'h047;
			{9'd302, 8'd129}: color_data = 12'h6df;
			{9'd302, 8'd130}: color_data = 12'heff;
			{9'd302, 8'd131}: color_data = 12'h6df;
			{9'd302, 8'd132}: color_data = 12'h0bf;
			{9'd302, 8'd133}: color_data = 12'h0be;
			{9'd302, 8'd134}: color_data = 12'h056;
			{9'd302, 8'd135}: color_data = 12'h012;
			{9'd302, 8'd136}: color_data = 12'h08b;
			{9'd302, 8'd137}: color_data = 12'h034;
			{9'd302, 8'd170}: color_data = 12'h000;
			{9'd302, 8'd171}: color_data = 12'h068;
			{9'd302, 8'd172}: color_data = 12'h8ef;
			{9'd302, 8'd173}: color_data = 12'hdff;
			{9'd302, 8'd174}: color_data = 12'h4cf;
			{9'd302, 8'd175}: color_data = 12'h0bf;
			{9'd302, 8'd176}: color_data = 12'h0ae;
			{9'd302, 8'd177}: color_data = 12'h035;
			{9'd302, 8'd178}: color_data = 12'h023;
			{9'd302, 8'd179}: color_data = 12'h08c;
			{9'd302, 8'd180}: color_data = 12'h023;
			{9'd302, 8'd204}: color_data = 12'h340;
			{9'd302, 8'd205}: color_data = 12'h9b0;
			{9'd302, 8'd206}: color_data = 12'hbc4;
			{9'd302, 8'd207}: color_data = 12'hfff;
			{9'd302, 8'd208}: color_data = 12'hefd;
			{9'd302, 8'd209}: color_data = 12'h9b1;
			{9'd302, 8'd210}: color_data = 12'h9b0;
			{9'd302, 8'd211}: color_data = 12'h9b0;
			{9'd302, 8'd212}: color_data = 12'h9b0;
			{9'd302, 8'd213}: color_data = 12'h9b0;
			{9'd302, 8'd214}: color_data = 12'h9b0;
			{9'd302, 8'd215}: color_data = 12'h780;
			{9'd302, 8'd216}: color_data = 12'h230;
			{9'd302, 8'd217}: color_data = 12'h020;
			{9'd302, 8'd218}: color_data = 12'h140;
			{9'd302, 8'd219}: color_data = 12'h350;
			{9'd302, 8'd220}: color_data = 12'h770;
			{9'd302, 8'd221}: color_data = 12'h440;
			{9'd302, 8'd222}: color_data = 12'h200;
			{9'd302, 8'd223}: color_data = 12'h900;
			{9'd302, 8'd224}: color_data = 12'hb00;
			{9'd302, 8'd225}: color_data = 12'h800;
			{9'd302, 8'd226}: color_data = 12'h200;
			{9'd302, 8'd227}: color_data = 12'hb30;
			{9'd302, 8'd228}: color_data = 12'hc10;
			{9'd302, 8'd229}: color_data = 12'h800;
			{9'd302, 8'd230}: color_data = 12'h300;
			{9'd302, 8'd231}: color_data = 12'h400;
			{9'd302, 8'd232}: color_data = 12'ha00;
			{9'd302, 8'd233}: color_data = 12'ha00;
			{9'd302, 8'd234}: color_data = 12'h500;
			{9'd302, 8'd235}: color_data = 12'h510;
			{9'd302, 8'd236}: color_data = 12'hd30;
			{9'd302, 8'd237}: color_data = 12'ha00;
			{9'd302, 8'd238}: color_data = 12'h700;
			{9'd302, 8'd239}: color_data = 12'h100;
			{9'd303, 8'd16}: color_data = 12'h010;
			{9'd303, 8'd17}: color_data = 12'h780;
			{9'd303, 8'd18}: color_data = 12'hac0;
			{9'd303, 8'd19}: color_data = 12'hdea;
			{9'd303, 8'd20}: color_data = 12'hfff;
			{9'd303, 8'd21}: color_data = 12'hcd7;
			{9'd303, 8'd22}: color_data = 12'h9b0;
			{9'd303, 8'd23}: color_data = 12'h9b0;
			{9'd303, 8'd24}: color_data = 12'h9b0;
			{9'd303, 8'd25}: color_data = 12'h9a0;
			{9'd303, 8'd26}: color_data = 12'h660;
			{9'd303, 8'd27}: color_data = 12'h130;
			{9'd303, 8'd28}: color_data = 12'h130;
			{9'd303, 8'd29}: color_data = 12'h240;
			{9'd303, 8'd30}: color_data = 12'h140;
			{9'd303, 8'd31}: color_data = 12'h240;
			{9'd303, 8'd32}: color_data = 12'h450;
			{9'd303, 8'd33}: color_data = 12'h460;
			{9'd303, 8'd34}: color_data = 12'h750;
			{9'd303, 8'd35}: color_data = 12'he10;
			{9'd303, 8'd36}: color_data = 12'he00;
			{9'd303, 8'd37}: color_data = 12'hb10;
			{9'd303, 8'd38}: color_data = 12'hd00;
			{9'd303, 8'd39}: color_data = 12'he00;
			{9'd303, 8'd40}: color_data = 12'hb10;
			{9'd303, 8'd41}: color_data = 12'hd00;
			{9'd303, 8'd42}: color_data = 12'hf00;
			{9'd303, 8'd43}: color_data = 12'h940;
			{9'd303, 8'd44}: color_data = 12'h450;
			{9'd303, 8'd45}: color_data = 12'h560;
			{9'd303, 8'd46}: color_data = 12'h8a0;
			{9'd303, 8'd47}: color_data = 12'h460;
			{9'd303, 8'd48}: color_data = 12'h140;
			{9'd303, 8'd49}: color_data = 12'h240;
			{9'd303, 8'd50}: color_data = 12'h020;
			{9'd303, 8'd51}: color_data = 12'h240;
			{9'd303, 8'd52}: color_data = 12'h560;
			{9'd303, 8'd53}: color_data = 12'h550;
			{9'd303, 8'd54}: color_data = 12'h550;
			{9'd303, 8'd55}: color_data = 12'h550;
			{9'd303, 8'd56}: color_data = 12'h550;
			{9'd303, 8'd57}: color_data = 12'h560;
			{9'd303, 8'd58}: color_data = 12'h760;
			{9'd303, 8'd59}: color_data = 12'h770;
			{9'd303, 8'd60}: color_data = 12'h660;
			{9'd303, 8'd61}: color_data = 12'h220;
			{9'd303, 8'd62}: color_data = 12'h000;
			{9'd303, 8'd68}: color_data = 12'h047;
			{9'd303, 8'd69}: color_data = 12'h6df;
			{9'd303, 8'd70}: color_data = 12'hfff;
			{9'd303, 8'd71}: color_data = 12'hdff;
			{9'd303, 8'd72}: color_data = 12'h5df;
			{9'd303, 8'd73}: color_data = 12'h068;
			{9'd303, 8'd74}: color_data = 12'h000;
			{9'd303, 8'd75}: color_data = 12'h012;
			{9'd303, 8'd76}: color_data = 12'h08c;
			{9'd303, 8'd77}: color_data = 12'h034;
			{9'd303, 8'd128}: color_data = 12'h047;
			{9'd303, 8'd129}: color_data = 12'h6df;
			{9'd303, 8'd130}: color_data = 12'hfff;
			{9'd303, 8'd131}: color_data = 12'hdff;
			{9'd303, 8'd132}: color_data = 12'h5df;
			{9'd303, 8'd133}: color_data = 12'h068;
			{9'd303, 8'd134}: color_data = 12'h000;
			{9'd303, 8'd135}: color_data = 12'h012;
			{9'd303, 8'd136}: color_data = 12'h08c;
			{9'd303, 8'd137}: color_data = 12'h034;
			{9'd303, 8'd170}: color_data = 12'h000;
			{9'd303, 8'd171}: color_data = 12'h068;
			{9'd303, 8'd172}: color_data = 12'h8ef;
			{9'd303, 8'd173}: color_data = 12'hfff;
			{9'd303, 8'd174}: color_data = 12'hcff;
			{9'd303, 8'd175}: color_data = 12'h4ce;
			{9'd303, 8'd176}: color_data = 12'h057;
			{9'd303, 8'd177}: color_data = 12'h000;
			{9'd303, 8'd178}: color_data = 12'h023;
			{9'd303, 8'd179}: color_data = 12'h08c;
			{9'd303, 8'd180}: color_data = 12'h023;
			{9'd303, 8'd204}: color_data = 12'h340;
			{9'd303, 8'd205}: color_data = 12'h9c0;
			{9'd303, 8'd206}: color_data = 12'hcd4;
			{9'd303, 8'd207}: color_data = 12'hfff;
			{9'd303, 8'd208}: color_data = 12'hffd;
			{9'd303, 8'd209}: color_data = 12'hac1;
			{9'd303, 8'd210}: color_data = 12'h9b0;
			{9'd303, 8'd211}: color_data = 12'hac0;
			{9'd303, 8'd212}: color_data = 12'hac0;
			{9'd303, 8'd213}: color_data = 12'hac0;
			{9'd303, 8'd214}: color_data = 12'hac0;
			{9'd303, 8'd215}: color_data = 12'h890;
			{9'd303, 8'd216}: color_data = 12'h230;
			{9'd303, 8'd217}: color_data = 12'h030;
			{9'd303, 8'd218}: color_data = 12'h140;
			{9'd303, 8'd219}: color_data = 12'h450;
			{9'd303, 8'd220}: color_data = 12'h770;
			{9'd303, 8'd221}: color_data = 12'h450;
			{9'd303, 8'd222}: color_data = 12'h200;
			{9'd303, 8'd223}: color_data = 12'h800;
			{9'd303, 8'd224}: color_data = 12'ha00;
			{9'd303, 8'd225}: color_data = 12'h700;
			{9'd303, 8'd226}: color_data = 12'h200;
			{9'd303, 8'd227}: color_data = 12'hb30;
			{9'd303, 8'd228}: color_data = 12'he20;
			{9'd303, 8'd229}: color_data = 12'ha00;
			{9'd303, 8'd230}: color_data = 12'h300;
			{9'd303, 8'd231}: color_data = 12'h400;
			{9'd303, 8'd232}: color_data = 12'ha00;
			{9'd303, 8'd233}: color_data = 12'ha00;
			{9'd303, 8'd234}: color_data = 12'h400;
			{9'd303, 8'd235}: color_data = 12'h510;
			{9'd303, 8'd236}: color_data = 12'hf40;
			{9'd303, 8'd237}: color_data = 12'hd10;
			{9'd303, 8'd238}: color_data = 12'h800;
			{9'd303, 8'd239}: color_data = 12'h100;
			{9'd304, 8'd16}: color_data = 12'h010;
			{9'd304, 8'd17}: color_data = 12'h780;
			{9'd304, 8'd18}: color_data = 12'hac0;
			{9'd304, 8'd19}: color_data = 12'hdea;
			{9'd304, 8'd20}: color_data = 12'hfff;
			{9'd304, 8'd21}: color_data = 12'hcd7;
			{9'd304, 8'd22}: color_data = 12'h8b0;
			{9'd304, 8'd23}: color_data = 12'h9b0;
			{9'd304, 8'd24}: color_data = 12'h9b0;
			{9'd304, 8'd25}: color_data = 12'h9b0;
			{9'd304, 8'd26}: color_data = 12'h9a0;
			{9'd304, 8'd27}: color_data = 12'h560;
			{9'd304, 8'd28}: color_data = 12'h120;
			{9'd304, 8'd29}: color_data = 12'h130;
			{9'd304, 8'd30}: color_data = 12'h240;
			{9'd304, 8'd31}: color_data = 12'h240;
			{9'd304, 8'd32}: color_data = 12'h140;
			{9'd304, 8'd33}: color_data = 12'h440;
			{9'd304, 8'd34}: color_data = 12'hc10;
			{9'd304, 8'd35}: color_data = 12'hf00;
			{9'd304, 8'd36}: color_data = 12'h720;
			{9'd304, 8'd37}: color_data = 12'h140;
			{9'd304, 8'd38}: color_data = 12'h920;
			{9'd304, 8'd39}: color_data = 12'hb10;
			{9'd304, 8'd40}: color_data = 12'h240;
			{9'd304, 8'd41}: color_data = 12'h530;
			{9'd304, 8'd42}: color_data = 12'he00;
			{9'd304, 8'd43}: color_data = 12'hd00;
			{9'd304, 8'd44}: color_data = 12'h430;
			{9'd304, 8'd45}: color_data = 12'h350;
			{9'd304, 8'd46}: color_data = 12'h790;
			{9'd304, 8'd47}: color_data = 12'h350;
			{9'd304, 8'd48}: color_data = 12'h030;
			{9'd304, 8'd49}: color_data = 12'h130;
			{9'd304, 8'd50}: color_data = 12'h020;
			{9'd304, 8'd51}: color_data = 12'h130;
			{9'd304, 8'd52}: color_data = 12'h240;
			{9'd304, 8'd53}: color_data = 12'h240;
			{9'd304, 8'd54}: color_data = 12'h240;
			{9'd304, 8'd55}: color_data = 12'h240;
			{9'd304, 8'd56}: color_data = 12'h240;
			{9'd304, 8'd57}: color_data = 12'h350;
			{9'd304, 8'd58}: color_data = 12'h560;
			{9'd304, 8'd59}: color_data = 12'h660;
			{9'd304, 8'd60}: color_data = 12'h760;
			{9'd304, 8'd61}: color_data = 12'h660;
			{9'd304, 8'd62}: color_data = 12'h220;
			{9'd304, 8'd63}: color_data = 12'h000;
			{9'd304, 8'd68}: color_data = 12'h047;
			{9'd304, 8'd69}: color_data = 12'h6df;
			{9'd304, 8'd70}: color_data = 12'hfff;
			{9'd304, 8'd71}: color_data = 12'hfff;
			{9'd304, 8'd72}: color_data = 12'h9aa;
			{9'd304, 8'd73}: color_data = 12'h011;
			{9'd304, 8'd75}: color_data = 12'h012;
			{9'd304, 8'd76}: color_data = 12'h08c;
			{9'd304, 8'd77}: color_data = 12'h034;
			{9'd304, 8'd128}: color_data = 12'h047;
			{9'd304, 8'd129}: color_data = 12'h6df;
			{9'd304, 8'd130}: color_data = 12'hfff;
			{9'd304, 8'd131}: color_data = 12'hfff;
			{9'd304, 8'd132}: color_data = 12'h9aa;
			{9'd304, 8'd133}: color_data = 12'h111;
			{9'd304, 8'd135}: color_data = 12'h012;
			{9'd304, 8'd136}: color_data = 12'h08c;
			{9'd304, 8'd137}: color_data = 12'h034;
			{9'd304, 8'd170}: color_data = 12'h000;
			{9'd304, 8'd171}: color_data = 12'h068;
			{9'd304, 8'd172}: color_data = 12'h7ef;
			{9'd304, 8'd173}: color_data = 12'hfff;
			{9'd304, 8'd174}: color_data = 12'hfff;
			{9'd304, 8'd175}: color_data = 12'h899;
			{9'd304, 8'd176}: color_data = 12'h001;
			{9'd304, 8'd178}: color_data = 12'h024;
			{9'd304, 8'd179}: color_data = 12'h08c;
			{9'd304, 8'd180}: color_data = 12'h023;
			{9'd304, 8'd204}: color_data = 12'h330;
			{9'd304, 8'd205}: color_data = 12'h790;
			{9'd304, 8'd206}: color_data = 12'h9b3;
			{9'd304, 8'd207}: color_data = 12'hcdd;
			{9'd304, 8'd208}: color_data = 12'hbca;
			{9'd304, 8'd209}: color_data = 12'h791;
			{9'd304, 8'd210}: color_data = 12'h790;
			{9'd304, 8'd211}: color_data = 12'h790;
			{9'd304, 8'd212}: color_data = 12'h790;
			{9'd304, 8'd213}: color_data = 12'h790;
			{9'd304, 8'd214}: color_data = 12'h790;
			{9'd304, 8'd215}: color_data = 12'h670;
			{9'd304, 8'd216}: color_data = 12'h230;
			{9'd304, 8'd217}: color_data = 12'h020;
			{9'd304, 8'd218}: color_data = 12'h130;
			{9'd304, 8'd219}: color_data = 12'h240;
			{9'd304, 8'd220}: color_data = 12'h550;
			{9'd304, 8'd221}: color_data = 12'h340;
			{9'd304, 8'd222}: color_data = 12'h200;
			{9'd304, 8'd223}: color_data = 12'h800;
			{9'd304, 8'd224}: color_data = 12'ha00;
			{9'd304, 8'd225}: color_data = 12'h800;
			{9'd304, 8'd226}: color_data = 12'h200;
			{9'd304, 8'd227}: color_data = 12'h920;
			{9'd304, 8'd228}: color_data = 12'hd30;
			{9'd304, 8'd229}: color_data = 12'h910;
			{9'd304, 8'd230}: color_data = 12'h200;
			{9'd304, 8'd231}: color_data = 12'h400;
			{9'd304, 8'd232}: color_data = 12'h900;
			{9'd304, 8'd233}: color_data = 12'ha00;
			{9'd304, 8'd234}: color_data = 12'h400;
			{9'd304, 8'd235}: color_data = 12'h310;
			{9'd304, 8'd236}: color_data = 12'hc30;
			{9'd304, 8'd237}: color_data = 12'hc20;
			{9'd304, 8'd238}: color_data = 12'h600;
			{9'd304, 8'd239}: color_data = 12'h000;
			{9'd305, 8'd16}: color_data = 12'h010;
			{9'd305, 8'd17}: color_data = 12'h780;
			{9'd305, 8'd18}: color_data = 12'hac0;
			{9'd305, 8'd19}: color_data = 12'hdea;
			{9'd305, 8'd20}: color_data = 12'hfff;
			{9'd305, 8'd21}: color_data = 12'hcd7;
			{9'd305, 8'd22}: color_data = 12'h9b0;
			{9'd305, 8'd23}: color_data = 12'h9b0;
			{9'd305, 8'd24}: color_data = 12'h9b0;
			{9'd305, 8'd25}: color_data = 12'h9b0;
			{9'd305, 8'd26}: color_data = 12'h9b0;
			{9'd305, 8'd27}: color_data = 12'h8a0;
			{9'd305, 8'd28}: color_data = 12'h450;
			{9'd305, 8'd29}: color_data = 12'h020;
			{9'd305, 8'd30}: color_data = 12'h130;
			{9'd305, 8'd31}: color_data = 12'h140;
			{9'd305, 8'd32}: color_data = 12'h140;
			{9'd305, 8'd33}: color_data = 12'ha10;
			{9'd305, 8'd34}: color_data = 12'hf00;
			{9'd305, 8'd35}: color_data = 12'h820;
			{9'd305, 8'd36}: color_data = 12'h140;
			{9'd305, 8'd37}: color_data = 12'h040;
			{9'd305, 8'd38}: color_data = 12'h820;
			{9'd305, 8'd39}: color_data = 12'ha10;
			{9'd305, 8'd40}: color_data = 12'h040;
			{9'd305, 8'd41}: color_data = 12'h040;
			{9'd305, 8'd42}: color_data = 12'h620;
			{9'd305, 8'd43}: color_data = 12'he00;
			{9'd305, 8'd44}: color_data = 12'hb00;
			{9'd305, 8'd45}: color_data = 12'h440;
			{9'd305, 8'd46}: color_data = 12'h7a0;
			{9'd305, 8'd47}: color_data = 12'h350;
			{9'd305, 8'd48}: color_data = 12'h010;
			{9'd305, 8'd49}: color_data = 12'h020;
			{9'd305, 8'd50}: color_data = 12'h020;
			{9'd305, 8'd51}: color_data = 12'h030;
			{9'd305, 8'd52}: color_data = 12'h140;
			{9'd305, 8'd53}: color_data = 12'h140;
			{9'd305, 8'd54}: color_data = 12'h140;
			{9'd305, 8'd55}: color_data = 12'h140;
			{9'd305, 8'd56}: color_data = 12'h140;
			{9'd305, 8'd57}: color_data = 12'h140;
			{9'd305, 8'd58}: color_data = 12'h240;
			{9'd305, 8'd59}: color_data = 12'h350;
			{9'd305, 8'd60}: color_data = 12'h660;
			{9'd305, 8'd61}: color_data = 12'h770;
			{9'd305, 8'd62}: color_data = 12'h550;
			{9'd305, 8'd63}: color_data = 12'h110;
			{9'd305, 8'd68}: color_data = 12'h047;
			{9'd305, 8'd69}: color_data = 12'h6df;
			{9'd305, 8'd70}: color_data = 12'hfff;
			{9'd305, 8'd71}: color_data = 12'hcbb;
			{9'd305, 8'd72}: color_data = 12'h323;
			{9'd305, 8'd73}: color_data = 12'h002;
			{9'd305, 8'd74}: color_data = 12'h000;
			{9'd305, 8'd75}: color_data = 12'h012;
			{9'd305, 8'd76}: color_data = 12'h08c;
			{9'd305, 8'd77}: color_data = 12'h034;
			{9'd305, 8'd128}: color_data = 12'h047;
			{9'd305, 8'd129}: color_data = 12'h6df;
			{9'd305, 8'd130}: color_data = 12'hfff;
			{9'd305, 8'd131}: color_data = 12'hcbb;
			{9'd305, 8'd132}: color_data = 12'h323;
			{9'd305, 8'd133}: color_data = 12'h002;
			{9'd305, 8'd134}: color_data = 12'h000;
			{9'd305, 8'd135}: color_data = 12'h012;
			{9'd305, 8'd136}: color_data = 12'h08c;
			{9'd305, 8'd137}: color_data = 12'h034;
			{9'd305, 8'd170}: color_data = 12'h000;
			{9'd305, 8'd171}: color_data = 12'h068;
			{9'd305, 8'd172}: color_data = 12'h8ef;
			{9'd305, 8'd173}: color_data = 12'hfff;
			{9'd305, 8'd174}: color_data = 12'haa9;
			{9'd305, 8'd175}: color_data = 12'h213;
			{9'd305, 8'd176}: color_data = 12'h002;
			{9'd305, 8'd178}: color_data = 12'h023;
			{9'd305, 8'd179}: color_data = 12'h08c;
			{9'd305, 8'd180}: color_data = 12'h023;
			{9'd305, 8'd204}: color_data = 12'h000;
			{9'd305, 8'd205}: color_data = 12'h120;
			{9'd305, 8'd206}: color_data = 12'h230;
			{9'd305, 8'd207}: color_data = 12'h242;
			{9'd305, 8'd208}: color_data = 12'h343;
			{9'd305, 8'd209}: color_data = 12'h241;
			{9'd305, 8'd210}: color_data = 12'h130;
			{9'd305, 8'd211}: color_data = 12'h130;
			{9'd305, 8'd212}: color_data = 12'h130;
			{9'd305, 8'd213}: color_data = 12'h130;
			{9'd305, 8'd214}: color_data = 12'h130;
			{9'd305, 8'd215}: color_data = 12'h130;
			{9'd305, 8'd216}: color_data = 12'h020;
			{9'd305, 8'd217}: color_data = 12'h020;
			{9'd305, 8'd218}: color_data = 12'h020;
			{9'd305, 8'd219}: color_data = 12'h020;
			{9'd305, 8'd220}: color_data = 12'h120;
			{9'd305, 8'd221}: color_data = 12'h000;
			{9'd305, 8'd222}: color_data = 12'h200;
			{9'd305, 8'd223}: color_data = 12'h900;
			{9'd305, 8'd224}: color_data = 12'ha00;
			{9'd305, 8'd225}: color_data = 12'h800;
			{9'd305, 8'd226}: color_data = 12'h100;
			{9'd305, 8'd227}: color_data = 12'h100;
			{9'd305, 8'd228}: color_data = 12'h310;
			{9'd305, 8'd229}: color_data = 12'h200;
			{9'd305, 8'd230}: color_data = 12'h000;
			{9'd305, 8'd231}: color_data = 12'h500;
			{9'd305, 8'd232}: color_data = 12'ha00;
			{9'd305, 8'd233}: color_data = 12'ha00;
			{9'd305, 8'd234}: color_data = 12'h500;
			{9'd305, 8'd235}: color_data = 12'h000;
			{9'd305, 8'd236}: color_data = 12'h200;
			{9'd305, 8'd237}: color_data = 12'h300;
			{9'd305, 8'd238}: color_data = 12'h100;
			{9'd305, 8'd239}: color_data = 12'h000;
			{9'd306, 8'd16}: color_data = 12'h010;
			{9'd306, 8'd17}: color_data = 12'h780;
			{9'd306, 8'd18}: color_data = 12'hac0;
			{9'd306, 8'd19}: color_data = 12'hdea;
			{9'd306, 8'd20}: color_data = 12'hfff;
			{9'd306, 8'd21}: color_data = 12'hffd;
			{9'd306, 8'd22}: color_data = 12'hbc5;
			{9'd306, 8'd23}: color_data = 12'h9b0;
			{9'd306, 8'd24}: color_data = 12'h9b0;
			{9'd306, 8'd25}: color_data = 12'h9b0;
			{9'd306, 8'd26}: color_data = 12'h9b0;
			{9'd306, 8'd27}: color_data = 12'h9b0;
			{9'd306, 8'd28}: color_data = 12'h890;
			{9'd306, 8'd29}: color_data = 12'h440;
			{9'd306, 8'd30}: color_data = 12'h020;
			{9'd306, 8'd31}: color_data = 12'h020;
			{9'd306, 8'd32}: color_data = 12'h120;
			{9'd306, 8'd33}: color_data = 12'hb00;
			{9'd306, 8'd34}: color_data = 12'h900;
			{9'd306, 8'd35}: color_data = 12'h120;
			{9'd306, 8'd36}: color_data = 12'h030;
			{9'd306, 8'd37}: color_data = 12'h020;
			{9'd306, 8'd38}: color_data = 12'h810;
			{9'd306, 8'd39}: color_data = 12'ha00;
			{9'd306, 8'd40}: color_data = 12'h020;
			{9'd306, 8'd41}: color_data = 12'h030;
			{9'd306, 8'd42}: color_data = 12'h020;
			{9'd306, 8'd43}: color_data = 12'h710;
			{9'd306, 8'd44}: color_data = 12'hc00;
			{9'd306, 8'd45}: color_data = 12'h431;
			{9'd306, 8'd46}: color_data = 12'hac8;
			{9'd306, 8'd47}: color_data = 12'h773;
			{9'd306, 8'd48}: color_data = 12'h340;
			{9'd306, 8'd49}: color_data = 12'h440;
			{9'd306, 8'd50}: color_data = 12'h130;
			{9'd306, 8'd51}: color_data = 12'h020;
			{9'd306, 8'd52}: color_data = 12'h020;
			{9'd306, 8'd53}: color_data = 12'h020;
			{9'd306, 8'd54}: color_data = 12'h020;
			{9'd306, 8'd55}: color_data = 12'h020;
			{9'd306, 8'd56}: color_data = 12'h020;
			{9'd306, 8'd57}: color_data = 12'h030;
			{9'd306, 8'd58}: color_data = 12'h140;
			{9'd306, 8'd59}: color_data = 12'h140;
			{9'd306, 8'd60}: color_data = 12'h350;
			{9'd306, 8'd61}: color_data = 12'h660;
			{9'd306, 8'd62}: color_data = 12'h770;
			{9'd306, 8'd63}: color_data = 12'h550;
			{9'd306, 8'd64}: color_data = 12'h110;
			{9'd306, 8'd68}: color_data = 12'h047;
			{9'd306, 8'd69}: color_data = 12'h6ef;
			{9'd306, 8'd70}: color_data = 12'hdcc;
			{9'd306, 8'd71}: color_data = 12'h434;
			{9'd306, 8'd72}: color_data = 12'h003;
			{9'd306, 8'd73}: color_data = 12'h005;
			{9'd306, 8'd74}: color_data = 12'h002;
			{9'd306, 8'd75}: color_data = 12'h012;
			{9'd306, 8'd76}: color_data = 12'h08c;
			{9'd306, 8'd77}: color_data = 12'h034;
			{9'd306, 8'd128}: color_data = 12'h047;
			{9'd306, 8'd129}: color_data = 12'h6ef;
			{9'd306, 8'd130}: color_data = 12'hddc;
			{9'd306, 8'd131}: color_data = 12'h434;
			{9'd306, 8'd132}: color_data = 12'h003;
			{9'd306, 8'd133}: color_data = 12'h005;
			{9'd306, 8'd134}: color_data = 12'h002;
			{9'd306, 8'd135}: color_data = 12'h012;
			{9'd306, 8'd136}: color_data = 12'h08c;
			{9'd306, 8'd137}: color_data = 12'h034;
			{9'd306, 8'd170}: color_data = 12'h000;
			{9'd306, 8'd171}: color_data = 12'h068;
			{9'd306, 8'd172}: color_data = 12'h8ff;
			{9'd306, 8'd173}: color_data = 12'hcbb;
			{9'd306, 8'd174}: color_data = 12'h223;
			{9'd306, 8'd175}: color_data = 12'h003;
			{9'd306, 8'd176}: color_data = 12'h005;
			{9'd306, 8'd177}: color_data = 12'h002;
			{9'd306, 8'd178}: color_data = 12'h023;
			{9'd306, 8'd179}: color_data = 12'h09c;
			{9'd306, 8'd180}: color_data = 12'h023;
			{9'd306, 8'd205}: color_data = 12'h110;
			{9'd306, 8'd206}: color_data = 12'h330;
			{9'd306, 8'd207}: color_data = 12'h452;
			{9'd306, 8'd208}: color_data = 12'h9a9;
			{9'd306, 8'd209}: color_data = 12'h9a9;
			{9'd306, 8'd210}: color_data = 12'h451;
			{9'd306, 8'd211}: color_data = 12'h330;
			{9'd306, 8'd212}: color_data = 12'h340;
			{9'd306, 8'd213}: color_data = 12'h340;
			{9'd306, 8'd214}: color_data = 12'h340;
			{9'd306, 8'd215}: color_data = 12'h120;
			{9'd306, 8'd216}: color_data = 12'h020;
			{9'd306, 8'd217}: color_data = 12'h130;
			{9'd306, 8'd218}: color_data = 12'h240;
			{9'd306, 8'd219}: color_data = 12'h450;
			{9'd306, 8'd220}: color_data = 12'h230;
			{9'd306, 8'd221}: color_data = 12'h000;
			{9'd306, 8'd222}: color_data = 12'h300;
			{9'd306, 8'd223}: color_data = 12'hc20;
			{9'd306, 8'd224}: color_data = 12'ha00;
			{9'd306, 8'd225}: color_data = 12'h800;
			{9'd306, 8'd226}: color_data = 12'h100;
			{9'd306, 8'd227}: color_data = 12'h300;
			{9'd306, 8'd228}: color_data = 12'h500;
			{9'd306, 8'd229}: color_data = 12'h500;
			{9'd306, 8'd230}: color_data = 12'h100;
			{9'd306, 8'd231}: color_data = 12'h710;
			{9'd306, 8'd232}: color_data = 12'hc10;
			{9'd306, 8'd233}: color_data = 12'h900;
			{9'd306, 8'd234}: color_data = 12'h500;
			{9'd306, 8'd235}: color_data = 12'h100;
			{9'd306, 8'd236}: color_data = 12'h500;
			{9'd306, 8'd237}: color_data = 12'h600;
			{9'd306, 8'd238}: color_data = 12'h400;
			{9'd306, 8'd239}: color_data = 12'h000;
			{9'd307, 8'd16}: color_data = 12'h010;
			{9'd307, 8'd17}: color_data = 12'h790;
			{9'd307, 8'd18}: color_data = 12'hac0;
			{9'd307, 8'd19}: color_data = 12'hbc5;
			{9'd307, 8'd20}: color_data = 12'hefd;
			{9'd307, 8'd21}: color_data = 12'hfff;
			{9'd307, 8'd22}: color_data = 12'hcd8;
			{9'd307, 8'd23}: color_data = 12'h8b0;
			{9'd307, 8'd24}: color_data = 12'h9b0;
			{9'd307, 8'd25}: color_data = 12'h9b0;
			{9'd307, 8'd26}: color_data = 12'h9b0;
			{9'd307, 8'd27}: color_data = 12'h9b0;
			{9'd307, 8'd28}: color_data = 12'h9b0;
			{9'd307, 8'd29}: color_data = 12'h780;
			{9'd307, 8'd30}: color_data = 12'h340;
			{9'd307, 8'd31}: color_data = 12'h230;
			{9'd307, 8'd32}: color_data = 12'h330;
			{9'd307, 8'd33}: color_data = 12'hc10;
			{9'd307, 8'd34}: color_data = 12'h730;
			{9'd307, 8'd35}: color_data = 12'h150;
			{9'd307, 8'd36}: color_data = 12'h240;
			{9'd307, 8'd37}: color_data = 12'h420;
			{9'd307, 8'd38}: color_data = 12'hc00;
			{9'd307, 8'd39}: color_data = 12'hd00;
			{9'd307, 8'd40}: color_data = 12'h620;
			{9'd307, 8'd41}: color_data = 12'h240;
			{9'd307, 8'd42}: color_data = 12'h150;
			{9'd307, 8'd43}: color_data = 12'h430;
			{9'd307, 8'd44}: color_data = 12'hc00;
			{9'd307, 8'd45}: color_data = 12'h742;
			{9'd307, 8'd46}: color_data = 12'hcdc;
			{9'd307, 8'd47}: color_data = 12'hbb4;
			{9'd307, 8'd48}: color_data = 12'h890;
			{9'd307, 8'd49}: color_data = 12'h890;
			{9'd307, 8'd50}: color_data = 12'h340;
			{9'd307, 8'd51}: color_data = 12'h120;
			{9'd307, 8'd52}: color_data = 12'h340;
			{9'd307, 8'd53}: color_data = 12'h230;
			{9'd307, 8'd54}: color_data = 12'h230;
			{9'd307, 8'd55}: color_data = 12'h230;
			{9'd307, 8'd56}: color_data = 12'h330;
			{9'd307, 8'd57}: color_data = 12'h230;
			{9'd307, 8'd58}: color_data = 12'h130;
			{9'd307, 8'd59}: color_data = 12'h140;
			{9'd307, 8'd60}: color_data = 12'h240;
			{9'd307, 8'd61}: color_data = 12'h350;
			{9'd307, 8'd62}: color_data = 12'h660;
			{9'd307, 8'd63}: color_data = 12'h760;
			{9'd307, 8'd64}: color_data = 12'h220;
			{9'd307, 8'd68}: color_data = 12'h057;
			{9'd307, 8'd69}: color_data = 12'h3bd;
			{9'd307, 8'd70}: color_data = 12'h555;
			{9'd307, 8'd71}: color_data = 12'h002;
			{9'd307, 8'd72}: color_data = 12'h005;
			{9'd307, 8'd73}: color_data = 12'h005;
			{9'd307, 8'd74}: color_data = 12'h004;
			{9'd307, 8'd75}: color_data = 12'h025;
			{9'd307, 8'd76}: color_data = 12'h09c;
			{9'd307, 8'd77}: color_data = 12'h034;
			{9'd307, 8'd128}: color_data = 12'h057;
			{9'd307, 8'd129}: color_data = 12'h3bd;
			{9'd307, 8'd130}: color_data = 12'h555;
			{9'd307, 8'd131}: color_data = 12'h002;
			{9'd307, 8'd132}: color_data = 12'h005;
			{9'd307, 8'd133}: color_data = 12'h005;
			{9'd307, 8'd134}: color_data = 12'h004;
			{9'd307, 8'd135}: color_data = 12'h024;
			{9'd307, 8'd136}: color_data = 12'h09c;
			{9'd307, 8'd137}: color_data = 12'h034;
			{9'd307, 8'd170}: color_data = 12'h000;
			{9'd307, 8'd171}: color_data = 12'h079;
			{9'd307, 8'd172}: color_data = 12'h4bd;
			{9'd307, 8'd173}: color_data = 12'h444;
			{9'd307, 8'd174}: color_data = 12'h002;
			{9'd307, 8'd175}: color_data = 12'h005;
			{9'd307, 8'd176}: color_data = 12'h005;
			{9'd307, 8'd177}: color_data = 12'h004;
			{9'd307, 8'd178}: color_data = 12'h036;
			{9'd307, 8'd179}: color_data = 12'h09c;
			{9'd307, 8'd180}: color_data = 12'h023;
			{9'd307, 8'd205}: color_data = 12'h230;
			{9'd307, 8'd206}: color_data = 12'h780;
			{9'd307, 8'd207}: color_data = 12'hab3;
			{9'd307, 8'd208}: color_data = 12'hfff;
			{9'd307, 8'd209}: color_data = 12'hffd;
			{9'd307, 8'd210}: color_data = 12'h9a2;
			{9'd307, 8'd211}: color_data = 12'h780;
			{9'd307, 8'd212}: color_data = 12'h890;
			{9'd307, 8'd213}: color_data = 12'h890;
			{9'd307, 8'd214}: color_data = 12'h770;
			{9'd307, 8'd215}: color_data = 12'h230;
			{9'd307, 8'd216}: color_data = 12'h030;
			{9'd307, 8'd217}: color_data = 12'h240;
			{9'd307, 8'd218}: color_data = 12'h450;
			{9'd307, 8'd219}: color_data = 12'h770;
			{9'd307, 8'd220}: color_data = 12'h440;
			{9'd307, 8'd221}: color_data = 12'h000;
			{9'd307, 8'd222}: color_data = 12'h410;
			{9'd307, 8'd223}: color_data = 12'hd30;
			{9'd307, 8'd224}: color_data = 12'hb00;
			{9'd307, 8'd225}: color_data = 12'h700;
			{9'd307, 8'd226}: color_data = 12'h200;
			{9'd307, 8'd227}: color_data = 12'h700;
			{9'd307, 8'd228}: color_data = 12'hb00;
			{9'd307, 8'd229}: color_data = 12'ha00;
			{9'd307, 8'd230}: color_data = 12'h300;
			{9'd307, 8'd231}: color_data = 12'h820;
			{9'd307, 8'd232}: color_data = 12'hd20;
			{9'd307, 8'd233}: color_data = 12'h900;
			{9'd307, 8'd234}: color_data = 12'h500;
			{9'd307, 8'd235}: color_data = 12'h300;
			{9'd307, 8'd236}: color_data = 12'h900;
			{9'd307, 8'd237}: color_data = 12'hb00;
			{9'd307, 8'd238}: color_data = 12'h800;
			{9'd307, 8'd239}: color_data = 12'h100;
			{9'd308, 8'd16}: color_data = 12'h000;
			{9'd308, 8'd17}: color_data = 12'h560;
			{9'd308, 8'd18}: color_data = 12'h8a0;
			{9'd308, 8'd19}: color_data = 12'h9b0;
			{9'd308, 8'd20}: color_data = 12'hdea;
			{9'd308, 8'd21}: color_data = 12'hfff;
			{9'd308, 8'd22}: color_data = 12'hdeb;
			{9'd308, 8'd23}: color_data = 12'hac2;
			{9'd308, 8'd24}: color_data = 12'h9b0;
			{9'd308, 8'd25}: color_data = 12'h9b0;
			{9'd308, 8'd26}: color_data = 12'h9b0;
			{9'd308, 8'd27}: color_data = 12'h9b0;
			{9'd308, 8'd28}: color_data = 12'h9b0;
			{9'd308, 8'd29}: color_data = 12'h9b0;
			{9'd308, 8'd30}: color_data = 12'h780;
			{9'd308, 8'd31}: color_data = 12'h780;
			{9'd308, 8'd32}: color_data = 12'h870;
			{9'd308, 8'd33}: color_data = 12'hd20;
			{9'd308, 8'd34}: color_data = 12'hc10;
			{9'd308, 8'd35}: color_data = 12'h940;
			{9'd308, 8'd36}: color_data = 12'ha40;
			{9'd308, 8'd37}: color_data = 12'hd10;
			{9'd308, 8'd38}: color_data = 12'hf33;
			{9'd308, 8'd39}: color_data = 12'hf34;
			{9'd308, 8'd40}: color_data = 12'he10;
			{9'd308, 8'd41}: color_data = 12'ha30;
			{9'd308, 8'd42}: color_data = 12'h940;
			{9'd308, 8'd43}: color_data = 12'hb20;
			{9'd308, 8'd44}: color_data = 12'hd00;
			{9'd308, 8'd45}: color_data = 12'h962;
			{9'd308, 8'd46}: color_data = 12'hdec;
			{9'd308, 8'd47}: color_data = 12'hbd4;
			{9'd308, 8'd48}: color_data = 12'h9b0;
			{9'd308, 8'd49}: color_data = 12'h9b0;
			{9'd308, 8'd50}: color_data = 12'h350;
			{9'd308, 8'd51}: color_data = 12'h330;
			{9'd308, 8'd52}: color_data = 12'h770;
			{9'd308, 8'd53}: color_data = 12'h780;
			{9'd308, 8'd54}: color_data = 12'h780;
			{9'd308, 8'd55}: color_data = 12'h780;
			{9'd308, 8'd56}: color_data = 12'h880;
			{9'd308, 8'd57}: color_data = 12'h670;
			{9'd308, 8'd58}: color_data = 12'h130;
			{9'd308, 8'd59}: color_data = 12'h030;
			{9'd308, 8'd60}: color_data = 12'h140;
			{9'd308, 8'd61}: color_data = 12'h240;
			{9'd308, 8'd62}: color_data = 12'h450;
			{9'd308, 8'd63}: color_data = 12'h660;
			{9'd308, 8'd64}: color_data = 12'h330;
			{9'd308, 8'd65}: color_data = 12'h000;
			{9'd308, 8'd68}: color_data = 12'h035;
			{9'd308, 8'd69}: color_data = 12'h047;
			{9'd308, 8'd70}: color_data = 12'h001;
			{9'd308, 8'd71}: color_data = 12'h004;
			{9'd308, 8'd72}: color_data = 12'h004;
			{9'd308, 8'd73}: color_data = 12'h004;
			{9'd308, 8'd74}: color_data = 12'h004;
			{9'd308, 8'd75}: color_data = 12'h015;
			{9'd308, 8'd76}: color_data = 12'h059;
			{9'd308, 8'd77}: color_data = 12'h023;
			{9'd308, 8'd128}: color_data = 12'h035;
			{9'd308, 8'd129}: color_data = 12'h047;
			{9'd308, 8'd130}: color_data = 12'h001;
			{9'd308, 8'd131}: color_data = 12'h004;
			{9'd308, 8'd132}: color_data = 12'h004;
			{9'd308, 8'd133}: color_data = 12'h004;
			{9'd308, 8'd134}: color_data = 12'h004;
			{9'd308, 8'd135}: color_data = 12'h015;
			{9'd308, 8'd136}: color_data = 12'h059;
			{9'd308, 8'd137}: color_data = 12'h023;
			{9'd308, 8'd170}: color_data = 12'h000;
			{9'd308, 8'd171}: color_data = 12'h047;
			{9'd308, 8'd172}: color_data = 12'h036;
			{9'd308, 8'd173}: color_data = 12'h001;
			{9'd308, 8'd174}: color_data = 12'h004;
			{9'd308, 8'd175}: color_data = 12'h004;
			{9'd308, 8'd176}: color_data = 12'h004;
			{9'd308, 8'd177}: color_data = 12'h004;
			{9'd308, 8'd178}: color_data = 12'h016;
			{9'd308, 8'd179}: color_data = 12'h059;
			{9'd308, 8'd180}: color_data = 12'h012;
			{9'd308, 8'd205}: color_data = 12'h330;
			{9'd308, 8'd206}: color_data = 12'h9b0;
			{9'd308, 8'd207}: color_data = 12'hbd3;
			{9'd308, 8'd208}: color_data = 12'hffe;
			{9'd308, 8'd209}: color_data = 12'hffd;
			{9'd308, 8'd210}: color_data = 12'hac2;
			{9'd308, 8'd211}: color_data = 12'h9b0;
			{9'd308, 8'd212}: color_data = 12'h9b0;
			{9'd308, 8'd213}: color_data = 12'h9b0;
			{9'd308, 8'd214}: color_data = 12'h780;
			{9'd308, 8'd215}: color_data = 12'h230;
			{9'd308, 8'd216}: color_data = 12'h030;
			{9'd308, 8'd217}: color_data = 12'h140;
			{9'd308, 8'd218}: color_data = 12'h450;
			{9'd308, 8'd219}: color_data = 12'h770;
			{9'd308, 8'd220}: color_data = 12'h440;
			{9'd308, 8'd221}: color_data = 12'h000;
			{9'd308, 8'd222}: color_data = 12'h410;
			{9'd308, 8'd223}: color_data = 12'he40;
			{9'd308, 8'd224}: color_data = 12'hd20;
			{9'd308, 8'd225}: color_data = 12'h800;
			{9'd308, 8'd226}: color_data = 12'h200;
			{9'd308, 8'd227}: color_data = 12'h600;
			{9'd308, 8'd228}: color_data = 12'ha00;
			{9'd308, 8'd229}: color_data = 12'h900;
			{9'd308, 8'd230}: color_data = 12'h300;
			{9'd308, 8'd231}: color_data = 12'h820;
			{9'd308, 8'd232}: color_data = 12'hf30;
			{9'd308, 8'd233}: color_data = 12'hc00;
			{9'd308, 8'd234}: color_data = 12'h500;
			{9'd308, 8'd235}: color_data = 12'h200;
			{9'd308, 8'd236}: color_data = 12'h900;
			{9'd308, 8'd237}: color_data = 12'ha00;
			{9'd308, 8'd238}: color_data = 12'h700;
			{9'd308, 8'd239}: color_data = 12'h100;
			{9'd309, 8'd17}: color_data = 12'h110;
			{9'd309, 8'd18}: color_data = 12'h780;
			{9'd309, 8'd19}: color_data = 12'hac0;
			{9'd309, 8'd20}: color_data = 12'hcd7;
			{9'd309, 8'd21}: color_data = 12'hfff;
			{9'd309, 8'd22}: color_data = 12'hfff;
			{9'd309, 8'd23}: color_data = 12'hde9;
			{9'd309, 8'd24}: color_data = 12'h9b1;
			{9'd309, 8'd25}: color_data = 12'h8b0;
			{9'd309, 8'd26}: color_data = 12'h9b0;
			{9'd309, 8'd27}: color_data = 12'h9b0;
			{9'd309, 8'd28}: color_data = 12'h9b0;
			{9'd309, 8'd29}: color_data = 12'h9b0;
			{9'd309, 8'd30}: color_data = 12'h9b0;
			{9'd309, 8'd31}: color_data = 12'h9b0;
			{9'd309, 8'd32}: color_data = 12'h9b0;
			{9'd309, 8'd33}: color_data = 12'he30;
			{9'd309, 8'd34}: color_data = 12'hf00;
			{9'd309, 8'd35}: color_data = 12'he10;
			{9'd309, 8'd36}: color_data = 12'he10;
			{9'd309, 8'd37}: color_data = 12'hf00;
			{9'd309, 8'd38}: color_data = 12'hf66;
			{9'd309, 8'd39}: color_data = 12'hf88;
			{9'd309, 8'd40}: color_data = 12'hf00;
			{9'd309, 8'd41}: color_data = 12'he10;
			{9'd309, 8'd42}: color_data = 12'he20;
			{9'd309, 8'd43}: color_data = 12'hf10;
			{9'd309, 8'd44}: color_data = 12'he00;
			{9'd309, 8'd45}: color_data = 12'h972;
			{9'd309, 8'd46}: color_data = 12'hdec;
			{9'd309, 8'd47}: color_data = 12'hbd4;
			{9'd309, 8'd48}: color_data = 12'h9b0;
			{9'd309, 8'd49}: color_data = 12'h9b0;
			{9'd309, 8'd50}: color_data = 12'h350;
			{9'd309, 8'd51}: color_data = 12'h330;
			{9'd309, 8'd52}: color_data = 12'h890;
			{9'd309, 8'd53}: color_data = 12'h9b0;
			{9'd309, 8'd54}: color_data = 12'h9b0;
			{9'd309, 8'd55}: color_data = 12'h9b0;
			{9'd309, 8'd56}: color_data = 12'h9b0;
			{9'd309, 8'd57}: color_data = 12'h9a0;
			{9'd309, 8'd58}: color_data = 12'h560;
			{9'd309, 8'd59}: color_data = 12'h130;
			{9'd309, 8'd60}: color_data = 12'h130;
			{9'd309, 8'd61}: color_data = 12'h140;
			{9'd309, 8'd62}: color_data = 12'h240;
			{9'd309, 8'd63}: color_data = 12'h560;
			{9'd309, 8'd64}: color_data = 12'h660;
			{9'd309, 8'd65}: color_data = 12'h220;
			{9'd309, 8'd68}: color_data = 12'h013;
			{9'd309, 8'd69}: color_data = 12'h027;
			{9'd309, 8'd70}: color_data = 12'h016;
			{9'd309, 8'd71}: color_data = 12'h027;
			{9'd309, 8'd72}: color_data = 12'h027;
			{9'd309, 8'd73}: color_data = 12'h027;
			{9'd309, 8'd74}: color_data = 12'h027;
			{9'd309, 8'd75}: color_data = 12'h028;
			{9'd309, 8'd76}: color_data = 12'h027;
			{9'd309, 8'd77}: color_data = 12'h001;
			{9'd309, 8'd128}: color_data = 12'h013;
			{9'd309, 8'd129}: color_data = 12'h027;
			{9'd309, 8'd130}: color_data = 12'h016;
			{9'd309, 8'd131}: color_data = 12'h027;
			{9'd309, 8'd132}: color_data = 12'h027;
			{9'd309, 8'd133}: color_data = 12'h027;
			{9'd309, 8'd134}: color_data = 12'h027;
			{9'd309, 8'd135}: color_data = 12'h028;
			{9'd309, 8'd136}: color_data = 12'h027;
			{9'd309, 8'd137}: color_data = 12'h001;
			{9'd309, 8'd170}: color_data = 12'h000;
			{9'd309, 8'd171}: color_data = 12'h014;
			{9'd309, 8'd172}: color_data = 12'h027;
			{9'd309, 8'd173}: color_data = 12'h016;
			{9'd309, 8'd174}: color_data = 12'h027;
			{9'd309, 8'd175}: color_data = 12'h027;
			{9'd309, 8'd176}: color_data = 12'h027;
			{9'd309, 8'd177}: color_data = 12'h027;
			{9'd309, 8'd178}: color_data = 12'h028;
			{9'd309, 8'd179}: color_data = 12'h026;
			{9'd309, 8'd180}: color_data = 12'h001;
			{9'd309, 8'd205}: color_data = 12'h330;
			{9'd309, 8'd206}: color_data = 12'h9b0;
			{9'd309, 8'd207}: color_data = 12'hbd3;
			{9'd309, 8'd208}: color_data = 12'hffe;
			{9'd309, 8'd209}: color_data = 12'hffd;
			{9'd309, 8'd210}: color_data = 12'hac2;
			{9'd309, 8'd211}: color_data = 12'h9b0;
			{9'd309, 8'd212}: color_data = 12'h9b0;
			{9'd309, 8'd213}: color_data = 12'h9b0;
			{9'd309, 8'd214}: color_data = 12'h780;
			{9'd309, 8'd215}: color_data = 12'h230;
			{9'd309, 8'd216}: color_data = 12'h030;
			{9'd309, 8'd217}: color_data = 12'h140;
			{9'd309, 8'd218}: color_data = 12'h450;
			{9'd309, 8'd219}: color_data = 12'h770;
			{9'd309, 8'd220}: color_data = 12'h440;
			{9'd309, 8'd221}: color_data = 12'h000;
			{9'd309, 8'd222}: color_data = 12'h200;
			{9'd309, 8'd223}: color_data = 12'hc30;
			{9'd309, 8'd224}: color_data = 12'hc30;
			{9'd309, 8'd225}: color_data = 12'h600;
			{9'd309, 8'd226}: color_data = 12'h100;
			{9'd309, 8'd227}: color_data = 12'h600;
			{9'd309, 8'd228}: color_data = 12'ha00;
			{9'd309, 8'd229}: color_data = 12'h900;
			{9'd309, 8'd230}: color_data = 12'h300;
			{9'd309, 8'd231}: color_data = 12'h620;
			{9'd309, 8'd232}: color_data = 12'hd40;
			{9'd309, 8'd233}: color_data = 12'ha20;
			{9'd309, 8'd234}: color_data = 12'h300;
			{9'd309, 8'd235}: color_data = 12'h200;
			{9'd309, 8'd236}: color_data = 12'h900;
			{9'd309, 8'd237}: color_data = 12'ha00;
			{9'd309, 8'd238}: color_data = 12'h700;
			{9'd309, 8'd239}: color_data = 12'h100;
			{9'd310, 8'd17}: color_data = 12'h000;
			{9'd310, 8'd18}: color_data = 12'h670;
			{9'd310, 8'd19}: color_data = 12'hac0;
			{9'd310, 8'd20}: color_data = 12'hac1;
			{9'd310, 8'd21}: color_data = 12'hde9;
			{9'd310, 8'd22}: color_data = 12'hfff;
			{9'd310, 8'd23}: color_data = 12'hfff;
			{9'd310, 8'd24}: color_data = 12'hcd8;
			{9'd310, 8'd25}: color_data = 12'h9b1;
			{9'd310, 8'd26}: color_data = 12'h9b0;
			{9'd310, 8'd27}: color_data = 12'h9b0;
			{9'd310, 8'd28}: color_data = 12'h9b0;
			{9'd310, 8'd29}: color_data = 12'h9b0;
			{9'd310, 8'd30}: color_data = 12'h9b0;
			{9'd310, 8'd31}: color_data = 12'h9c0;
			{9'd310, 8'd32}: color_data = 12'h9b0;
			{9'd310, 8'd33}: color_data = 12'he30;
			{9'd310, 8'd34}: color_data = 12'hc50;
			{9'd310, 8'd35}: color_data = 12'h870;
			{9'd310, 8'd36}: color_data = 12'h970;
			{9'd310, 8'd37}: color_data = 12'hd50;
			{9'd310, 8'd38}: color_data = 12'hf11;
			{9'd310, 8'd39}: color_data = 12'hf22;
			{9'd310, 8'd40}: color_data = 12'hd10;
			{9'd310, 8'd41}: color_data = 12'h960;
			{9'd310, 8'd42}: color_data = 12'haa0;
			{9'd310, 8'd43}: color_data = 12'hc70;
			{9'd310, 8'd44}: color_data = 12'he20;
			{9'd310, 8'd45}: color_data = 12'hb92;
			{9'd310, 8'd46}: color_data = 12'hdfc;
			{9'd310, 8'd47}: color_data = 12'hbc4;
			{9'd310, 8'd48}: color_data = 12'h9b0;
			{9'd310, 8'd49}: color_data = 12'h9b0;
			{9'd310, 8'd50}: color_data = 12'h350;
			{9'd310, 8'd51}: color_data = 12'h230;
			{9'd310, 8'd52}: color_data = 12'h890;
			{9'd310, 8'd53}: color_data = 12'h9c0;
			{9'd310, 8'd54}: color_data = 12'h9b0;
			{9'd310, 8'd55}: color_data = 12'h9b0;
			{9'd310, 8'd56}: color_data = 12'h9b0;
			{9'd310, 8'd57}: color_data = 12'h9b0;
			{9'd310, 8'd58}: color_data = 12'h8a0;
			{9'd310, 8'd59}: color_data = 12'h550;
			{9'd310, 8'd60}: color_data = 12'h120;
			{9'd310, 8'd61}: color_data = 12'h130;
			{9'd310, 8'd62}: color_data = 12'h240;
			{9'd310, 8'd63}: color_data = 12'h560;
			{9'd310, 8'd64}: color_data = 12'h770;
			{9'd310, 8'd65}: color_data = 12'h220;
			{9'd310, 8'd68}: color_data = 12'h046;
			{9'd310, 8'd69}: color_data = 12'h09e;
			{9'd310, 8'd70}: color_data = 12'h09e;
			{9'd310, 8'd71}: color_data = 12'h09e;
			{9'd310, 8'd72}: color_data = 12'h09e;
			{9'd310, 8'd73}: color_data = 12'h09e;
			{9'd310, 8'd74}: color_data = 12'h09e;
			{9'd310, 8'd75}: color_data = 12'h09e;
			{9'd310, 8'd76}: color_data = 12'h08c;
			{9'd310, 8'd77}: color_data = 12'h023;
			{9'd310, 8'd128}: color_data = 12'h045;
			{9'd310, 8'd129}: color_data = 12'h09e;
			{9'd310, 8'd130}: color_data = 12'h0ae;
			{9'd310, 8'd131}: color_data = 12'h09e;
			{9'd310, 8'd132}: color_data = 12'h09e;
			{9'd310, 8'd133}: color_data = 12'h09e;
			{9'd310, 8'd134}: color_data = 12'h09e;
			{9'd310, 8'd135}: color_data = 12'h09e;
			{9'd310, 8'd136}: color_data = 12'h08c;
			{9'd310, 8'd137}: color_data = 12'h023;
			{9'd310, 8'd170}: color_data = 12'h000;
			{9'd310, 8'd171}: color_data = 12'h057;
			{9'd310, 8'd172}: color_data = 12'h0ae;
			{9'd310, 8'd173}: color_data = 12'h09e;
			{9'd310, 8'd174}: color_data = 12'h09e;
			{9'd310, 8'd175}: color_data = 12'h09e;
			{9'd310, 8'd176}: color_data = 12'h09e;
			{9'd310, 8'd177}: color_data = 12'h09e;
			{9'd310, 8'd178}: color_data = 12'h09e;
			{9'd310, 8'd179}: color_data = 12'h07b;
			{9'd310, 8'd180}: color_data = 12'h012;
			{9'd310, 8'd205}: color_data = 12'h330;
			{9'd310, 8'd206}: color_data = 12'h9b0;
			{9'd310, 8'd207}: color_data = 12'hbc3;
			{9'd310, 8'd208}: color_data = 12'hffe;
			{9'd310, 8'd209}: color_data = 12'hffd;
			{9'd310, 8'd210}: color_data = 12'hac2;
			{9'd310, 8'd211}: color_data = 12'h9b0;
			{9'd310, 8'd212}: color_data = 12'h9b0;
			{9'd310, 8'd213}: color_data = 12'h9b0;
			{9'd310, 8'd214}: color_data = 12'h780;
			{9'd310, 8'd215}: color_data = 12'h230;
			{9'd310, 8'd216}: color_data = 12'h030;
			{9'd310, 8'd217}: color_data = 12'h140;
			{9'd310, 8'd218}: color_data = 12'h450;
			{9'd310, 8'd219}: color_data = 12'h770;
			{9'd310, 8'd220}: color_data = 12'h440;
			{9'd310, 8'd221}: color_data = 12'h000;
			{9'd310, 8'd222}: color_data = 12'h000;
			{9'd310, 8'd223}: color_data = 12'h200;
			{9'd310, 8'd224}: color_data = 12'h300;
			{9'd310, 8'd225}: color_data = 12'h100;
			{9'd310, 8'd226}: color_data = 12'h000;
			{9'd310, 8'd227}: color_data = 12'h700;
			{9'd310, 8'd228}: color_data = 12'ha00;
			{9'd310, 8'd229}: color_data = 12'h900;
			{9'd310, 8'd230}: color_data = 12'h300;
			{9'd310, 8'd231}: color_data = 12'h100;
			{9'd310, 8'd232}: color_data = 12'h310;
			{9'd310, 8'd233}: color_data = 12'h200;
			{9'd310, 8'd234}: color_data = 12'h000;
			{9'd310, 8'd235}: color_data = 12'h300;
			{9'd310, 8'd236}: color_data = 12'h900;
			{9'd310, 8'd237}: color_data = 12'ha00;
			{9'd310, 8'd238}: color_data = 12'h700;
			{9'd310, 8'd239}: color_data = 12'h100;
			{9'd311, 8'd18}: color_data = 12'h220;
			{9'd311, 8'd19}: color_data = 12'h790;
			{9'd311, 8'd20}: color_data = 12'h9c0;
			{9'd311, 8'd21}: color_data = 12'hac2;
			{9'd311, 8'd22}: color_data = 12'hdea;
			{9'd311, 8'd23}: color_data = 12'hfff;
			{9'd311, 8'd24}: color_data = 12'hffe;
			{9'd311, 8'd25}: color_data = 12'heeb;
			{9'd311, 8'd26}: color_data = 12'hcd7;
			{9'd311, 8'd27}: color_data = 12'h9b0;
			{9'd311, 8'd28}: color_data = 12'h9b0;
			{9'd311, 8'd29}: color_data = 12'h9b0;
			{9'd311, 8'd30}: color_data = 12'h9b0;
			{9'd311, 8'd31}: color_data = 12'h9b0;
			{9'd311, 8'd32}: color_data = 12'h9a0;
			{9'd311, 8'd33}: color_data = 12'he30;
			{9'd311, 8'd34}: color_data = 12'hb70;
			{9'd311, 8'd35}: color_data = 12'h690;
			{9'd311, 8'd36}: color_data = 12'h7a0;
			{9'd311, 8'd37}: color_data = 12'haa0;
			{9'd311, 8'd38}: color_data = 12'he30;
			{9'd311, 8'd39}: color_data = 12'he20;
			{9'd311, 8'd40}: color_data = 12'h970;
			{9'd311, 8'd41}: color_data = 12'h680;
			{9'd311, 8'd42}: color_data = 12'h8d0;
			{9'd311, 8'd43}: color_data = 12'haa0;
			{9'd311, 8'd44}: color_data = 12'he20;
			{9'd311, 8'd45}: color_data = 12'hba2;
			{9'd311, 8'd46}: color_data = 12'hefc;
			{9'd311, 8'd47}: color_data = 12'hbc4;
			{9'd311, 8'd48}: color_data = 12'h9b0;
			{9'd311, 8'd49}: color_data = 12'h9b0;
			{9'd311, 8'd50}: color_data = 12'h350;
			{9'd311, 8'd51}: color_data = 12'h230;
			{9'd311, 8'd52}: color_data = 12'h880;
			{9'd311, 8'd53}: color_data = 12'h9b0;
			{9'd311, 8'd54}: color_data = 12'h9b0;
			{9'd311, 8'd55}: color_data = 12'h9b0;
			{9'd311, 8'd56}: color_data = 12'h9b0;
			{9'd311, 8'd57}: color_data = 12'h9b0;
			{9'd311, 8'd58}: color_data = 12'h9b0;
			{9'd311, 8'd59}: color_data = 12'h660;
			{9'd311, 8'd60}: color_data = 12'h020;
			{9'd311, 8'd61}: color_data = 12'h130;
			{9'd311, 8'd62}: color_data = 12'h240;
			{9'd311, 8'd63}: color_data = 12'h560;
			{9'd311, 8'd64}: color_data = 12'h760;
			{9'd311, 8'd65}: color_data = 12'h220;
			{9'd311, 8'd68}: color_data = 12'h057;
			{9'd311, 8'd69}: color_data = 12'h4ef;
			{9'd311, 8'd70}: color_data = 12'h7ef;
			{9'd311, 8'd71}: color_data = 12'h0cf;
			{9'd311, 8'd72}: color_data = 12'h0cf;
			{9'd311, 8'd73}: color_data = 12'h0df;
			{9'd311, 8'd74}: color_data = 12'h0bd;
			{9'd311, 8'd75}: color_data = 12'h068;
			{9'd311, 8'd76}: color_data = 12'h09c;
			{9'd311, 8'd77}: color_data = 12'h034;
			{9'd311, 8'd128}: color_data = 12'h057;
			{9'd311, 8'd129}: color_data = 12'h4ef;
			{9'd311, 8'd130}: color_data = 12'h7ef;
			{9'd311, 8'd131}: color_data = 12'h0cf;
			{9'd311, 8'd132}: color_data = 12'h0cf;
			{9'd311, 8'd133}: color_data = 12'h0df;
			{9'd311, 8'd134}: color_data = 12'h0bd;
			{9'd311, 8'd135}: color_data = 12'h068;
			{9'd311, 8'd136}: color_data = 12'h09c;
			{9'd311, 8'd137}: color_data = 12'h034;
			{9'd311, 8'd170}: color_data = 12'h000;
			{9'd311, 8'd171}: color_data = 12'h069;
			{9'd311, 8'd172}: color_data = 12'h6ef;
			{9'd311, 8'd173}: color_data = 12'h6ef;
			{9'd311, 8'd174}: color_data = 12'h0cf;
			{9'd311, 8'd175}: color_data = 12'h0cf;
			{9'd311, 8'd176}: color_data = 12'h0df;
			{9'd311, 8'd177}: color_data = 12'h0ac;
			{9'd311, 8'd178}: color_data = 12'h079;
			{9'd311, 8'd179}: color_data = 12'h09c;
			{9'd311, 8'd180}: color_data = 12'h023;
			{9'd311, 8'd205}: color_data = 12'h330;
			{9'd311, 8'd206}: color_data = 12'h9b0;
			{9'd311, 8'd207}: color_data = 12'hbc3;
			{9'd311, 8'd208}: color_data = 12'hffe;
			{9'd311, 8'd209}: color_data = 12'hffd;
			{9'd311, 8'd210}: color_data = 12'hac2;
			{9'd311, 8'd211}: color_data = 12'h9b0;
			{9'd311, 8'd212}: color_data = 12'h9b0;
			{9'd311, 8'd213}: color_data = 12'h9b0;
			{9'd311, 8'd214}: color_data = 12'h780;
			{9'd311, 8'd215}: color_data = 12'h230;
			{9'd311, 8'd216}: color_data = 12'h030;
			{9'd311, 8'd217}: color_data = 12'h140;
			{9'd311, 8'd218}: color_data = 12'h450;
			{9'd311, 8'd219}: color_data = 12'h770;
			{9'd311, 8'd220}: color_data = 12'h440;
			{9'd311, 8'd221}: color_data = 12'h000;
			{9'd311, 8'd222}: color_data = 12'h100;
			{9'd311, 8'd223}: color_data = 12'h500;
			{9'd311, 8'd224}: color_data = 12'h600;
			{9'd311, 8'd225}: color_data = 12'h400;
			{9'd311, 8'd226}: color_data = 12'h100;
			{9'd311, 8'd227}: color_data = 12'ha20;
			{9'd311, 8'd228}: color_data = 12'hb10;
			{9'd311, 8'd229}: color_data = 12'h900;
			{9'd311, 8'd230}: color_data = 12'h300;
			{9'd311, 8'd231}: color_data = 12'h200;
			{9'd311, 8'd232}: color_data = 12'h500;
			{9'd311, 8'd233}: color_data = 12'h500;
			{9'd311, 8'd234}: color_data = 12'h200;
			{9'd311, 8'd235}: color_data = 12'h410;
			{9'd311, 8'd236}: color_data = 12'hc20;
			{9'd311, 8'd237}: color_data = 12'ha00;
			{9'd311, 8'd238}: color_data = 12'h700;
			{9'd311, 8'd239}: color_data = 12'h100;
			{9'd312, 8'd19}: color_data = 12'h230;
			{9'd312, 8'd20}: color_data = 12'h8a0;
			{9'd312, 8'd21}: color_data = 12'h9c0;
			{9'd312, 8'd22}: color_data = 12'hac3;
			{9'd312, 8'd23}: color_data = 12'heec;
			{9'd312, 8'd24}: color_data = 12'hfff;
			{9'd312, 8'd25}: color_data = 12'hfff;
			{9'd312, 8'd26}: color_data = 12'hffe;
			{9'd312, 8'd27}: color_data = 12'hbd6;
			{9'd312, 8'd28}: color_data = 12'hab1;
			{9'd312, 8'd29}: color_data = 12'hcd7;
			{9'd312, 8'd30}: color_data = 12'hcd7;
			{9'd312, 8'd31}: color_data = 12'h9c1;
			{9'd312, 8'd32}: color_data = 12'h9a0;
			{9'd312, 8'd33}: color_data = 12'he20;
			{9'd312, 8'd34}: color_data = 12'he20;
			{9'd312, 8'd35}: color_data = 12'h980;
			{9'd312, 8'd36}: color_data = 12'h790;
			{9'd312, 8'd37}: color_data = 12'h8b0;
			{9'd312, 8'd38}: color_data = 12'hc60;
			{9'd312, 8'd39}: color_data = 12'hd40;
			{9'd312, 8'd40}: color_data = 12'h8a0;
			{9'd312, 8'd41}: color_data = 12'h680;
			{9'd312, 8'd42}: color_data = 12'h9a0;
			{9'd312, 8'd43}: color_data = 12'hd40;
			{9'd312, 8'd44}: color_data = 12'he00;
			{9'd312, 8'd45}: color_data = 12'ha82;
			{9'd312, 8'd46}: color_data = 12'hdec;
			{9'd312, 8'd47}: color_data = 12'hbc4;
			{9'd312, 8'd48}: color_data = 12'h8b0;
			{9'd312, 8'd49}: color_data = 12'h8b0;
			{9'd312, 8'd50}: color_data = 12'h350;
			{9'd312, 8'd51}: color_data = 12'h564;
			{9'd312, 8'd52}: color_data = 12'hcd9;
			{9'd312, 8'd53}: color_data = 12'hbc4;
			{9'd312, 8'd54}: color_data = 12'h9b0;
			{9'd312, 8'd55}: color_data = 12'h9b0;
			{9'd312, 8'd56}: color_data = 12'h9b0;
			{9'd312, 8'd57}: color_data = 12'h9b0;
			{9'd312, 8'd58}: color_data = 12'h9a0;
			{9'd312, 8'd59}: color_data = 12'h560;
			{9'd312, 8'd60}: color_data = 12'h020;
			{9'd312, 8'd61}: color_data = 12'h130;
			{9'd312, 8'd62}: color_data = 12'h240;
			{9'd312, 8'd63}: color_data = 12'h560;
			{9'd312, 8'd64}: color_data = 12'h760;
			{9'd312, 8'd65}: color_data = 12'h220;
			{9'd312, 8'd68}: color_data = 12'h047;
			{9'd312, 8'd69}: color_data = 12'h6df;
			{9'd312, 8'd70}: color_data = 12'heff;
			{9'd312, 8'd71}: color_data = 12'h6df;
			{9'd312, 8'd72}: color_data = 12'h0bf;
			{9'd312, 8'd73}: color_data = 12'h0bf;
			{9'd312, 8'd74}: color_data = 12'h056;
			{9'd312, 8'd75}: color_data = 12'h012;
			{9'd312, 8'd76}: color_data = 12'h08b;
			{9'd312, 8'd77}: color_data = 12'h034;
			{9'd312, 8'd128}: color_data = 12'h047;
			{9'd312, 8'd129}: color_data = 12'h6df;
			{9'd312, 8'd130}: color_data = 12'heff;
			{9'd312, 8'd131}: color_data = 12'h6df;
			{9'd312, 8'd132}: color_data = 12'h0bf;
			{9'd312, 8'd133}: color_data = 12'h0bf;
			{9'd312, 8'd134}: color_data = 12'h056;
			{9'd312, 8'd135}: color_data = 12'h012;
			{9'd312, 8'd136}: color_data = 12'h08b;
			{9'd312, 8'd137}: color_data = 12'h034;
			{9'd312, 8'd170}: color_data = 12'h000;
			{9'd312, 8'd171}: color_data = 12'h068;
			{9'd312, 8'd172}: color_data = 12'h8ef;
			{9'd312, 8'd173}: color_data = 12'hdff;
			{9'd312, 8'd174}: color_data = 12'h4cf;
			{9'd312, 8'd175}: color_data = 12'h0bf;
			{9'd312, 8'd176}: color_data = 12'h0ae;
			{9'd312, 8'd177}: color_data = 12'h035;
			{9'd312, 8'd178}: color_data = 12'h023;
			{9'd312, 8'd179}: color_data = 12'h08c;
			{9'd312, 8'd180}: color_data = 12'h023;
			{9'd312, 8'd205}: color_data = 12'h330;
			{9'd312, 8'd206}: color_data = 12'h9b0;
			{9'd312, 8'd207}: color_data = 12'hbc3;
			{9'd312, 8'd208}: color_data = 12'hffe;
			{9'd312, 8'd209}: color_data = 12'hffd;
			{9'd312, 8'd210}: color_data = 12'hac2;
			{9'd312, 8'd211}: color_data = 12'h9b0;
			{9'd312, 8'd212}: color_data = 12'h9b0;
			{9'd312, 8'd213}: color_data = 12'h9b0;
			{9'd312, 8'd214}: color_data = 12'h780;
			{9'd312, 8'd215}: color_data = 12'h230;
			{9'd312, 8'd216}: color_data = 12'h030;
			{9'd312, 8'd217}: color_data = 12'h140;
			{9'd312, 8'd218}: color_data = 12'h450;
			{9'd312, 8'd219}: color_data = 12'h770;
			{9'd312, 8'd220}: color_data = 12'h440;
			{9'd312, 8'd221}: color_data = 12'h000;
			{9'd312, 8'd222}: color_data = 12'h200;
			{9'd312, 8'd223}: color_data = 12'h900;
			{9'd312, 8'd224}: color_data = 12'hb00;
			{9'd312, 8'd225}: color_data = 12'h800;
			{9'd312, 8'd226}: color_data = 12'h200;
			{9'd312, 8'd227}: color_data = 12'hb30;
			{9'd312, 8'd228}: color_data = 12'hc10;
			{9'd312, 8'd229}: color_data = 12'h800;
			{9'd312, 8'd230}: color_data = 12'h300;
			{9'd312, 8'd231}: color_data = 12'h400;
			{9'd312, 8'd232}: color_data = 12'ha00;
			{9'd312, 8'd233}: color_data = 12'ha00;
			{9'd312, 8'd234}: color_data = 12'h500;
			{9'd312, 8'd235}: color_data = 12'h510;
			{9'd312, 8'd236}: color_data = 12'hd30;
			{9'd312, 8'd237}: color_data = 12'ha00;
			{9'd312, 8'd238}: color_data = 12'h700;
			{9'd312, 8'd239}: color_data = 12'h100;
			{9'd313, 8'd19}: color_data = 12'h000;
			{9'd313, 8'd20}: color_data = 12'h340;
			{9'd313, 8'd21}: color_data = 12'h8a0;
			{9'd313, 8'd22}: color_data = 12'h9b0;
			{9'd313, 8'd23}: color_data = 12'hbc4;
			{9'd313, 8'd24}: color_data = 12'hdea;
			{9'd313, 8'd25}: color_data = 12'hefc;
			{9'd313, 8'd26}: color_data = 12'hfff;
			{9'd313, 8'd27}: color_data = 12'heeb;
			{9'd313, 8'd28}: color_data = 12'hac3;
			{9'd313, 8'd29}: color_data = 12'hffd;
			{9'd313, 8'd30}: color_data = 12'hffe;
			{9'd313, 8'd31}: color_data = 12'hac3;
			{9'd313, 8'd32}: color_data = 12'h9b0;
			{9'd313, 8'd33}: color_data = 12'hc50;
			{9'd313, 8'd34}: color_data = 12'hf00;
			{9'd313, 8'd35}: color_data = 12'hd40;
			{9'd313, 8'd36}: color_data = 12'h880;
			{9'd313, 8'd37}: color_data = 12'h6a0;
			{9'd313, 8'd38}: color_data = 12'hb50;
			{9'd313, 8'd39}: color_data = 12'hd30;
			{9'd313, 8'd40}: color_data = 12'h690;
			{9'd313, 8'd41}: color_data = 12'h680;
			{9'd313, 8'd42}: color_data = 12'hc50;
			{9'd313, 8'd43}: color_data = 12'hf00;
			{9'd313, 8'd44}: color_data = 12'hc10;
			{9'd313, 8'd45}: color_data = 12'h882;
			{9'd313, 8'd46}: color_data = 12'hdec;
			{9'd313, 8'd47}: color_data = 12'hde8;
			{9'd313, 8'd48}: color_data = 12'hbd4;
			{9'd313, 8'd49}: color_data = 12'hbc5;
			{9'd313, 8'd50}: color_data = 12'h351;
			{9'd313, 8'd51}: color_data = 12'h898;
			{9'd313, 8'd52}: color_data = 12'hfff;
			{9'd313, 8'd53}: color_data = 12'heeb;
			{9'd313, 8'd54}: color_data = 12'hac2;
			{9'd313, 8'd55}: color_data = 12'h9b0;
			{9'd313, 8'd56}: color_data = 12'h9b0;
			{9'd313, 8'd57}: color_data = 12'h9b0;
			{9'd313, 8'd58}: color_data = 12'h9a0;
			{9'd313, 8'd59}: color_data = 12'h560;
			{9'd313, 8'd60}: color_data = 12'h020;
			{9'd313, 8'd61}: color_data = 12'h130;
			{9'd313, 8'd62}: color_data = 12'h240;
			{9'd313, 8'd63}: color_data = 12'h560;
			{9'd313, 8'd64}: color_data = 12'h760;
			{9'd313, 8'd65}: color_data = 12'h220;
			{9'd313, 8'd68}: color_data = 12'h047;
			{9'd313, 8'd69}: color_data = 12'h6df;
			{9'd313, 8'd70}: color_data = 12'hfff;
			{9'd313, 8'd71}: color_data = 12'hdff;
			{9'd313, 8'd72}: color_data = 12'h5df;
			{9'd313, 8'd73}: color_data = 12'h068;
			{9'd313, 8'd74}: color_data = 12'h000;
			{9'd313, 8'd75}: color_data = 12'h012;
			{9'd313, 8'd76}: color_data = 12'h08c;
			{9'd313, 8'd77}: color_data = 12'h034;
			{9'd313, 8'd128}: color_data = 12'h047;
			{9'd313, 8'd129}: color_data = 12'h6df;
			{9'd313, 8'd130}: color_data = 12'hfff;
			{9'd313, 8'd131}: color_data = 12'hdff;
			{9'd313, 8'd132}: color_data = 12'h5df;
			{9'd313, 8'd133}: color_data = 12'h068;
			{9'd313, 8'd134}: color_data = 12'h000;
			{9'd313, 8'd135}: color_data = 12'h012;
			{9'd313, 8'd136}: color_data = 12'h08c;
			{9'd313, 8'd137}: color_data = 12'h034;
			{9'd313, 8'd170}: color_data = 12'h000;
			{9'd313, 8'd171}: color_data = 12'h068;
			{9'd313, 8'd172}: color_data = 12'h8ef;
			{9'd313, 8'd173}: color_data = 12'hfff;
			{9'd313, 8'd174}: color_data = 12'hcff;
			{9'd313, 8'd175}: color_data = 12'h4ce;
			{9'd313, 8'd176}: color_data = 12'h057;
			{9'd313, 8'd177}: color_data = 12'h000;
			{9'd313, 8'd178}: color_data = 12'h023;
			{9'd313, 8'd179}: color_data = 12'h08c;
			{9'd313, 8'd180}: color_data = 12'h023;
			{9'd313, 8'd205}: color_data = 12'h330;
			{9'd313, 8'd206}: color_data = 12'h9b0;
			{9'd313, 8'd207}: color_data = 12'hbc3;
			{9'd313, 8'd208}: color_data = 12'hffe;
			{9'd313, 8'd209}: color_data = 12'hffd;
			{9'd313, 8'd210}: color_data = 12'hac2;
			{9'd313, 8'd211}: color_data = 12'h9b0;
			{9'd313, 8'd212}: color_data = 12'h9b0;
			{9'd313, 8'd213}: color_data = 12'h9b0;
			{9'd313, 8'd214}: color_data = 12'h780;
			{9'd313, 8'd215}: color_data = 12'h230;
			{9'd313, 8'd216}: color_data = 12'h030;
			{9'd313, 8'd217}: color_data = 12'h140;
			{9'd313, 8'd218}: color_data = 12'h450;
			{9'd313, 8'd219}: color_data = 12'h770;
			{9'd313, 8'd220}: color_data = 12'h440;
			{9'd313, 8'd221}: color_data = 12'h000;
			{9'd313, 8'd222}: color_data = 12'h200;
			{9'd313, 8'd223}: color_data = 12'h900;
			{9'd313, 8'd224}: color_data = 12'ha00;
			{9'd313, 8'd225}: color_data = 12'h700;
			{9'd313, 8'd226}: color_data = 12'h200;
			{9'd313, 8'd227}: color_data = 12'hb30;
			{9'd313, 8'd228}: color_data = 12'he20;
			{9'd313, 8'd229}: color_data = 12'ha00;
			{9'd313, 8'd230}: color_data = 12'h300;
			{9'd313, 8'd231}: color_data = 12'h400;
			{9'd313, 8'd232}: color_data = 12'ha00;
			{9'd313, 8'd233}: color_data = 12'ha00;
			{9'd313, 8'd234}: color_data = 12'h400;
			{9'd313, 8'd235}: color_data = 12'h510;
			{9'd313, 8'd236}: color_data = 12'hf40;
			{9'd313, 8'd237}: color_data = 12'hd10;
			{9'd313, 8'd238}: color_data = 12'h800;
			{9'd313, 8'd239}: color_data = 12'h100;
			{9'd314, 8'd20}: color_data = 12'h000;
			{9'd314, 8'd21}: color_data = 12'h450;
			{9'd314, 8'd22}: color_data = 12'h9b0;
			{9'd314, 8'd23}: color_data = 12'hac0;
			{9'd314, 8'd24}: color_data = 12'h9b0;
			{9'd314, 8'd25}: color_data = 12'hbc5;
			{9'd314, 8'd26}: color_data = 12'hefd;
			{9'd314, 8'd27}: color_data = 12'hde9;
			{9'd314, 8'd28}: color_data = 12'hac3;
			{9'd314, 8'd29}: color_data = 12'heeb;
			{9'd314, 8'd30}: color_data = 12'heec;
			{9'd314, 8'd31}: color_data = 12'hac2;
			{9'd314, 8'd32}: color_data = 12'h8b0;
			{9'd314, 8'd33}: color_data = 12'h9b0;
			{9'd314, 8'd34}: color_data = 12'hd40;
			{9'd314, 8'd35}: color_data = 12'hf00;
			{9'd314, 8'd36}: color_data = 12'hd50;
			{9'd314, 8'd37}: color_data = 12'h870;
			{9'd314, 8'd38}: color_data = 12'hc20;
			{9'd314, 8'd39}: color_data = 12'hd10;
			{9'd314, 8'd40}: color_data = 12'h750;
			{9'd314, 8'd41}: color_data = 12'ha30;
			{9'd314, 8'd42}: color_data = 12'hf00;
			{9'd314, 8'd43}: color_data = 12'hd20;
			{9'd314, 8'd44}: color_data = 12'h760;
			{9'd314, 8'd45}: color_data = 12'h9b1;
			{9'd314, 8'd46}: color_data = 12'hefc;
			{9'd314, 8'd47}: color_data = 12'hfff;
			{9'd314, 8'd48}: color_data = 12'hfff;
			{9'd314, 8'd49}: color_data = 12'hffe;
			{9'd314, 8'd50}: color_data = 12'h565;
			{9'd314, 8'd51}: color_data = 12'h786;
			{9'd314, 8'd52}: color_data = 12'hfff;
			{9'd314, 8'd53}: color_data = 12'hfff;
			{9'd314, 8'd54}: color_data = 12'hdea;
			{9'd314, 8'd55}: color_data = 12'hab1;
			{9'd314, 8'd56}: color_data = 12'h9b0;
			{9'd314, 8'd57}: color_data = 12'h9b0;
			{9'd314, 8'd58}: color_data = 12'h9a0;
			{9'd314, 8'd59}: color_data = 12'h560;
			{9'd314, 8'd60}: color_data = 12'h020;
			{9'd314, 8'd61}: color_data = 12'h130;
			{9'd314, 8'd62}: color_data = 12'h240;
			{9'd314, 8'd63}: color_data = 12'h560;
			{9'd314, 8'd64}: color_data = 12'h760;
			{9'd314, 8'd65}: color_data = 12'h220;
			{9'd314, 8'd68}: color_data = 12'h047;
			{9'd314, 8'd69}: color_data = 12'h6df;
			{9'd314, 8'd70}: color_data = 12'hfff;
			{9'd314, 8'd71}: color_data = 12'hfff;
			{9'd314, 8'd72}: color_data = 12'h9aa;
			{9'd314, 8'd73}: color_data = 12'h011;
			{9'd314, 8'd75}: color_data = 12'h012;
			{9'd314, 8'd76}: color_data = 12'h08c;
			{9'd314, 8'd77}: color_data = 12'h034;
			{9'd314, 8'd128}: color_data = 12'h047;
			{9'd314, 8'd129}: color_data = 12'h6df;
			{9'd314, 8'd130}: color_data = 12'hfff;
			{9'd314, 8'd131}: color_data = 12'hfff;
			{9'd314, 8'd132}: color_data = 12'h9aa;
			{9'd314, 8'd133}: color_data = 12'h111;
			{9'd314, 8'd135}: color_data = 12'h012;
			{9'd314, 8'd136}: color_data = 12'h08c;
			{9'd314, 8'd137}: color_data = 12'h034;
			{9'd314, 8'd170}: color_data = 12'h000;
			{9'd314, 8'd171}: color_data = 12'h068;
			{9'd314, 8'd172}: color_data = 12'h7ef;
			{9'd314, 8'd173}: color_data = 12'hfff;
			{9'd314, 8'd174}: color_data = 12'hfff;
			{9'd314, 8'd175}: color_data = 12'h899;
			{9'd314, 8'd176}: color_data = 12'h001;
			{9'd314, 8'd178}: color_data = 12'h024;
			{9'd314, 8'd179}: color_data = 12'h08c;
			{9'd314, 8'd180}: color_data = 12'h023;
			{9'd314, 8'd205}: color_data = 12'h330;
			{9'd314, 8'd206}: color_data = 12'h9b0;
			{9'd314, 8'd207}: color_data = 12'hbc3;
			{9'd314, 8'd208}: color_data = 12'hffe;
			{9'd314, 8'd209}: color_data = 12'hffd;
			{9'd314, 8'd210}: color_data = 12'hac2;
			{9'd314, 8'd211}: color_data = 12'h9b0;
			{9'd314, 8'd212}: color_data = 12'h9b0;
			{9'd314, 8'd213}: color_data = 12'h9b0;
			{9'd314, 8'd214}: color_data = 12'h780;
			{9'd314, 8'd215}: color_data = 12'h230;
			{9'd314, 8'd216}: color_data = 12'h030;
			{9'd314, 8'd217}: color_data = 12'h140;
			{9'd314, 8'd218}: color_data = 12'h450;
			{9'd314, 8'd219}: color_data = 12'h770;
			{9'd314, 8'd220}: color_data = 12'h440;
			{9'd314, 8'd221}: color_data = 12'h000;
			{9'd314, 8'd222}: color_data = 12'h200;
			{9'd314, 8'd223}: color_data = 12'h800;
			{9'd314, 8'd224}: color_data = 12'ha00;
			{9'd314, 8'd225}: color_data = 12'h800;
			{9'd314, 8'd226}: color_data = 12'h200;
			{9'd314, 8'd227}: color_data = 12'h930;
			{9'd314, 8'd228}: color_data = 12'hd30;
			{9'd314, 8'd229}: color_data = 12'h910;
			{9'd314, 8'd230}: color_data = 12'h200;
			{9'd314, 8'd231}: color_data = 12'h400;
			{9'd314, 8'd232}: color_data = 12'h900;
			{9'd314, 8'd233}: color_data = 12'ha00;
			{9'd314, 8'd234}: color_data = 12'h400;
			{9'd314, 8'd235}: color_data = 12'h310;
			{9'd314, 8'd236}: color_data = 12'hc30;
			{9'd314, 8'd237}: color_data = 12'hc20;
			{9'd314, 8'd238}: color_data = 12'h600;
			{9'd314, 8'd239}: color_data = 12'h000;
			{9'd315, 8'd21}: color_data = 12'h000;
			{9'd315, 8'd22}: color_data = 12'h560;
			{9'd315, 8'd23}: color_data = 12'h9b0;
			{9'd315, 8'd24}: color_data = 12'h8b0;
			{9'd315, 8'd25}: color_data = 12'h9b0;
			{9'd315, 8'd26}: color_data = 12'hac3;
			{9'd315, 8'd27}: color_data = 12'hac2;
			{9'd315, 8'd28}: color_data = 12'h9c0;
			{9'd315, 8'd29}: color_data = 12'hac2;
			{9'd315, 8'd30}: color_data = 12'hac2;
			{9'd315, 8'd31}: color_data = 12'h9b0;
			{9'd315, 8'd32}: color_data = 12'h9b0;
			{9'd315, 8'd33}: color_data = 12'h9c0;
			{9'd315, 8'd34}: color_data = 12'hab0;
			{9'd315, 8'd35}: color_data = 12'he40;
			{9'd315, 8'd36}: color_data = 12'hf10;
			{9'd315, 8'd37}: color_data = 12'he20;
			{9'd315, 8'd38}: color_data = 12'hf10;
			{9'd315, 8'd39}: color_data = 12'hf10;
			{9'd315, 8'd40}: color_data = 12'he10;
			{9'd315, 8'd41}: color_data = 12'hf10;
			{9'd315, 8'd42}: color_data = 12'he20;
			{9'd315, 8'd43}: color_data = 12'ha90;
			{9'd315, 8'd44}: color_data = 12'h8b0;
			{9'd315, 8'd45}: color_data = 12'hac1;
			{9'd315, 8'd46}: color_data = 12'hefc;
			{9'd315, 8'd47}: color_data = 12'hfff;
			{9'd315, 8'd48}: color_data = 12'hfff;
			{9'd315, 8'd49}: color_data = 12'hffe;
			{9'd315, 8'd50}: color_data = 12'h565;
			{9'd315, 8'd51}: color_data = 12'h460;
			{9'd315, 8'd52}: color_data = 12'hde8;
			{9'd315, 8'd53}: color_data = 12'hfff;
			{9'd315, 8'd54}: color_data = 12'hfff;
			{9'd315, 8'd55}: color_data = 12'hdd8;
			{9'd315, 8'd56}: color_data = 12'h9b0;
			{9'd315, 8'd57}: color_data = 12'h9b0;
			{9'd315, 8'd58}: color_data = 12'h9a0;
			{9'd315, 8'd59}: color_data = 12'h560;
			{9'd315, 8'd60}: color_data = 12'h020;
			{9'd315, 8'd61}: color_data = 12'h130;
			{9'd315, 8'd62}: color_data = 12'h240;
			{9'd315, 8'd63}: color_data = 12'h560;
			{9'd315, 8'd64}: color_data = 12'h760;
			{9'd315, 8'd65}: color_data = 12'h220;
			{9'd315, 8'd68}: color_data = 12'h047;
			{9'd315, 8'd69}: color_data = 12'h6df;
			{9'd315, 8'd70}: color_data = 12'hfff;
			{9'd315, 8'd71}: color_data = 12'hcbb;
			{9'd315, 8'd72}: color_data = 12'h323;
			{9'd315, 8'd73}: color_data = 12'h002;
			{9'd315, 8'd74}: color_data = 12'h000;
			{9'd315, 8'd75}: color_data = 12'h012;
			{9'd315, 8'd76}: color_data = 12'h08c;
			{9'd315, 8'd77}: color_data = 12'h034;
			{9'd315, 8'd128}: color_data = 12'h047;
			{9'd315, 8'd129}: color_data = 12'h6df;
			{9'd315, 8'd130}: color_data = 12'hfff;
			{9'd315, 8'd131}: color_data = 12'hcbb;
			{9'd315, 8'd132}: color_data = 12'h323;
			{9'd315, 8'd133}: color_data = 12'h002;
			{9'd315, 8'd134}: color_data = 12'h000;
			{9'd315, 8'd135}: color_data = 12'h012;
			{9'd315, 8'd136}: color_data = 12'h08c;
			{9'd315, 8'd137}: color_data = 12'h034;
			{9'd315, 8'd170}: color_data = 12'h000;
			{9'd315, 8'd171}: color_data = 12'h068;
			{9'd315, 8'd172}: color_data = 12'h8ef;
			{9'd315, 8'd173}: color_data = 12'hfff;
			{9'd315, 8'd174}: color_data = 12'haa9;
			{9'd315, 8'd175}: color_data = 12'h213;
			{9'd315, 8'd176}: color_data = 12'h002;
			{9'd315, 8'd178}: color_data = 12'h023;
			{9'd315, 8'd179}: color_data = 12'h08c;
			{9'd315, 8'd180}: color_data = 12'h023;
			{9'd315, 8'd205}: color_data = 12'h330;
			{9'd315, 8'd206}: color_data = 12'h9b0;
			{9'd315, 8'd207}: color_data = 12'hbc3;
			{9'd315, 8'd208}: color_data = 12'hffe;
			{9'd315, 8'd209}: color_data = 12'hffd;
			{9'd315, 8'd210}: color_data = 12'hac2;
			{9'd315, 8'd211}: color_data = 12'h9b0;
			{9'd315, 8'd212}: color_data = 12'h9b0;
			{9'd315, 8'd213}: color_data = 12'h9b0;
			{9'd315, 8'd214}: color_data = 12'h780;
			{9'd315, 8'd215}: color_data = 12'h230;
			{9'd315, 8'd216}: color_data = 12'h030;
			{9'd315, 8'd217}: color_data = 12'h140;
			{9'd315, 8'd218}: color_data = 12'h450;
			{9'd315, 8'd219}: color_data = 12'h770;
			{9'd315, 8'd220}: color_data = 12'h440;
			{9'd315, 8'd221}: color_data = 12'h000;
			{9'd315, 8'd222}: color_data = 12'h200;
			{9'd315, 8'd223}: color_data = 12'h900;
			{9'd315, 8'd224}: color_data = 12'ha00;
			{9'd315, 8'd225}: color_data = 12'h800;
			{9'd315, 8'd226}: color_data = 12'h100;
			{9'd315, 8'd227}: color_data = 12'h100;
			{9'd315, 8'd228}: color_data = 12'h310;
			{9'd315, 8'd229}: color_data = 12'h200;
			{9'd315, 8'd230}: color_data = 12'h000;
			{9'd315, 8'd231}: color_data = 12'h500;
			{9'd315, 8'd232}: color_data = 12'ha00;
			{9'd315, 8'd233}: color_data = 12'ha00;
			{9'd315, 8'd234}: color_data = 12'h500;
			{9'd315, 8'd235}: color_data = 12'h000;
			{9'd315, 8'd236}: color_data = 12'h200;
			{9'd315, 8'd237}: color_data = 12'h300;
			{9'd315, 8'd238}: color_data = 12'h100;
			{9'd315, 8'd239}: color_data = 12'h000;
			{9'd316, 8'd22}: color_data = 12'h110;
			{9'd316, 8'd23}: color_data = 12'h230;
			{9'd316, 8'd24}: color_data = 12'h560;
			{9'd316, 8'd25}: color_data = 12'h9c0;
			{9'd316, 8'd26}: color_data = 12'h9b0;
			{9'd316, 8'd27}: color_data = 12'h9b0;
			{9'd316, 8'd28}: color_data = 12'h9b0;
			{9'd316, 8'd29}: color_data = 12'h9b0;
			{9'd316, 8'd30}: color_data = 12'h9b0;
			{9'd316, 8'd31}: color_data = 12'h9b0;
			{9'd316, 8'd32}: color_data = 12'h9b0;
			{9'd316, 8'd33}: color_data = 12'h9c0;
			{9'd316, 8'd34}: color_data = 12'h9c0;
			{9'd316, 8'd35}: color_data = 12'haa0;
			{9'd316, 8'd36}: color_data = 12'hc70;
			{9'd316, 8'd37}: color_data = 12'hc70;
			{9'd316, 8'd38}: color_data = 12'hc80;
			{9'd316, 8'd39}: color_data = 12'hc80;
			{9'd316, 8'd40}: color_data = 12'hc70;
			{9'd316, 8'd41}: color_data = 12'hc70;
			{9'd316, 8'd42}: color_data = 12'hb90;
			{9'd316, 8'd43}: color_data = 12'h9c0;
			{9'd316, 8'd44}: color_data = 12'h9c0;
			{9'd316, 8'd45}: color_data = 12'hac2;
			{9'd316, 8'd46}: color_data = 12'hefc;
			{9'd316, 8'd47}: color_data = 12'hdd8;
			{9'd316, 8'd48}: color_data = 12'hbd4;
			{9'd316, 8'd49}: color_data = 12'hbd5;
			{9'd316, 8'd50}: color_data = 12'h461;
			{9'd316, 8'd51}: color_data = 12'h460;
			{9'd316, 8'd52}: color_data = 12'hac1;
			{9'd316, 8'd53}: color_data = 12'hdea;
			{9'd316, 8'd54}: color_data = 12'hfff;
			{9'd316, 8'd55}: color_data = 12'hdea;
			{9'd316, 8'd56}: color_data = 12'h9b0;
			{9'd316, 8'd57}: color_data = 12'h9b0;
			{9'd316, 8'd58}: color_data = 12'h9a0;
			{9'd316, 8'd59}: color_data = 12'h560;
			{9'd316, 8'd60}: color_data = 12'h020;
			{9'd316, 8'd61}: color_data = 12'h130;
			{9'd316, 8'd62}: color_data = 12'h240;
			{9'd316, 8'd63}: color_data = 12'h560;
			{9'd316, 8'd64}: color_data = 12'h760;
			{9'd316, 8'd65}: color_data = 12'h220;
			{9'd316, 8'd68}: color_data = 12'h047;
			{9'd316, 8'd69}: color_data = 12'h6ef;
			{9'd316, 8'd70}: color_data = 12'hddc;
			{9'd316, 8'd71}: color_data = 12'h434;
			{9'd316, 8'd72}: color_data = 12'h003;
			{9'd316, 8'd73}: color_data = 12'h005;
			{9'd316, 8'd74}: color_data = 12'h002;
			{9'd316, 8'd75}: color_data = 12'h012;
			{9'd316, 8'd76}: color_data = 12'h08c;
			{9'd316, 8'd77}: color_data = 12'h034;
			{9'd316, 8'd128}: color_data = 12'h047;
			{9'd316, 8'd129}: color_data = 12'h6ef;
			{9'd316, 8'd130}: color_data = 12'hddc;
			{9'd316, 8'd131}: color_data = 12'h434;
			{9'd316, 8'd132}: color_data = 12'h003;
			{9'd316, 8'd133}: color_data = 12'h005;
			{9'd316, 8'd134}: color_data = 12'h002;
			{9'd316, 8'd135}: color_data = 12'h012;
			{9'd316, 8'd136}: color_data = 12'h08c;
			{9'd316, 8'd137}: color_data = 12'h034;
			{9'd316, 8'd170}: color_data = 12'h000;
			{9'd316, 8'd171}: color_data = 12'h068;
			{9'd316, 8'd172}: color_data = 12'h8ff;
			{9'd316, 8'd173}: color_data = 12'hcbb;
			{9'd316, 8'd174}: color_data = 12'h323;
			{9'd316, 8'd175}: color_data = 12'h003;
			{9'd316, 8'd176}: color_data = 12'h005;
			{9'd316, 8'd177}: color_data = 12'h002;
			{9'd316, 8'd178}: color_data = 12'h023;
			{9'd316, 8'd179}: color_data = 12'h09c;
			{9'd316, 8'd180}: color_data = 12'h023;
			{9'd316, 8'd205}: color_data = 12'h330;
			{9'd316, 8'd206}: color_data = 12'h9b0;
			{9'd316, 8'd207}: color_data = 12'hbc3;
			{9'd316, 8'd208}: color_data = 12'hffe;
			{9'd316, 8'd209}: color_data = 12'hffd;
			{9'd316, 8'd210}: color_data = 12'hac2;
			{9'd316, 8'd211}: color_data = 12'h9b0;
			{9'd316, 8'd212}: color_data = 12'h9b0;
			{9'd316, 8'd213}: color_data = 12'h9b0;
			{9'd316, 8'd214}: color_data = 12'h780;
			{9'd316, 8'd215}: color_data = 12'h230;
			{9'd316, 8'd216}: color_data = 12'h030;
			{9'd316, 8'd217}: color_data = 12'h140;
			{9'd316, 8'd218}: color_data = 12'h450;
			{9'd316, 8'd219}: color_data = 12'h770;
			{9'd316, 8'd220}: color_data = 12'h440;
			{9'd316, 8'd221}: color_data = 12'h000;
			{9'd316, 8'd222}: color_data = 12'h300;
			{9'd316, 8'd223}: color_data = 12'hc20;
			{9'd316, 8'd224}: color_data = 12'ha00;
			{9'd316, 8'd225}: color_data = 12'h800;
			{9'd316, 8'd226}: color_data = 12'h100;
			{9'd316, 8'd227}: color_data = 12'h300;
			{9'd316, 8'd228}: color_data = 12'h500;
			{9'd316, 8'd229}: color_data = 12'h500;
			{9'd316, 8'd230}: color_data = 12'h100;
			{9'd316, 8'd231}: color_data = 12'h710;
			{9'd316, 8'd232}: color_data = 12'hc10;
			{9'd316, 8'd233}: color_data = 12'h900;
			{9'd316, 8'd234}: color_data = 12'h500;
			{9'd316, 8'd235}: color_data = 12'h100;
			{9'd316, 8'd236}: color_data = 12'h500;
			{9'd316, 8'd237}: color_data = 12'h600;
			{9'd316, 8'd238}: color_data = 12'h400;
			{9'd316, 8'd239}: color_data = 12'h000;
			{9'd317, 8'd24}: color_data = 12'h120;
			{9'd317, 8'd25}: color_data = 12'h450;
			{9'd317, 8'd26}: color_data = 12'h450;
			{9'd317, 8'd27}: color_data = 12'h450;
			{9'd317, 8'd28}: color_data = 12'h450;
			{9'd317, 8'd29}: color_data = 12'h450;
			{9'd317, 8'd30}: color_data = 12'h450;
			{9'd317, 8'd31}: color_data = 12'h450;
			{9'd317, 8'd32}: color_data = 12'h450;
			{9'd317, 8'd33}: color_data = 12'h450;
			{9'd317, 8'd34}: color_data = 12'h450;
			{9'd317, 8'd35}: color_data = 12'h460;
			{9'd317, 8'd36}: color_data = 12'h460;
			{9'd317, 8'd37}: color_data = 12'h460;
			{9'd317, 8'd38}: color_data = 12'h460;
			{9'd317, 8'd39}: color_data = 12'h460;
			{9'd317, 8'd40}: color_data = 12'h460;
			{9'd317, 8'd41}: color_data = 12'h460;
			{9'd317, 8'd42}: color_data = 12'h460;
			{9'd317, 8'd43}: color_data = 12'h450;
			{9'd317, 8'd44}: color_data = 12'h450;
			{9'd317, 8'd45}: color_data = 12'h662;
			{9'd317, 8'd46}: color_data = 12'hdec;
			{9'd317, 8'd47}: color_data = 12'hbd4;
			{9'd317, 8'd48}: color_data = 12'h9c0;
			{9'd317, 8'd49}: color_data = 12'h9c0;
			{9'd317, 8'd50}: color_data = 12'h340;
			{9'd317, 8'd51}: color_data = 12'h460;
			{9'd317, 8'd52}: color_data = 12'h9b0;
			{9'd317, 8'd53}: color_data = 12'hcd7;
			{9'd317, 8'd54}: color_data = 12'hfff;
			{9'd317, 8'd55}: color_data = 12'hdea;
			{9'd317, 8'd56}: color_data = 12'h9b0;
			{9'd317, 8'd57}: color_data = 12'h9b0;
			{9'd317, 8'd58}: color_data = 12'h9a0;
			{9'd317, 8'd59}: color_data = 12'h560;
			{9'd317, 8'd60}: color_data = 12'h020;
			{9'd317, 8'd61}: color_data = 12'h130;
			{9'd317, 8'd62}: color_data = 12'h240;
			{9'd317, 8'd63}: color_data = 12'h560;
			{9'd317, 8'd64}: color_data = 12'h760;
			{9'd317, 8'd65}: color_data = 12'h220;
			{9'd317, 8'd68}: color_data = 12'h057;
			{9'd317, 8'd69}: color_data = 12'h3bd;
			{9'd317, 8'd70}: color_data = 12'h555;
			{9'd317, 8'd71}: color_data = 12'h002;
			{9'd317, 8'd72}: color_data = 12'h005;
			{9'd317, 8'd73}: color_data = 12'h005;
			{9'd317, 8'd74}: color_data = 12'h004;
			{9'd317, 8'd75}: color_data = 12'h025;
			{9'd317, 8'd76}: color_data = 12'h09c;
			{9'd317, 8'd77}: color_data = 12'h034;
			{9'd317, 8'd128}: color_data = 12'h057;
			{9'd317, 8'd129}: color_data = 12'h3bd;
			{9'd317, 8'd130}: color_data = 12'h555;
			{9'd317, 8'd131}: color_data = 12'h002;
			{9'd317, 8'd132}: color_data = 12'h005;
			{9'd317, 8'd133}: color_data = 12'h005;
			{9'd317, 8'd134}: color_data = 12'h004;
			{9'd317, 8'd135}: color_data = 12'h025;
			{9'd317, 8'd136}: color_data = 12'h09c;
			{9'd317, 8'd137}: color_data = 12'h034;
			{9'd317, 8'd170}: color_data = 12'h000;
			{9'd317, 8'd171}: color_data = 12'h079;
			{9'd317, 8'd172}: color_data = 12'h4bd;
			{9'd317, 8'd173}: color_data = 12'h444;
			{9'd317, 8'd174}: color_data = 12'h002;
			{9'd317, 8'd175}: color_data = 12'h005;
			{9'd317, 8'd176}: color_data = 12'h005;
			{9'd317, 8'd177}: color_data = 12'h004;
			{9'd317, 8'd178}: color_data = 12'h036;
			{9'd317, 8'd179}: color_data = 12'h09c;
			{9'd317, 8'd180}: color_data = 12'h023;
			{9'd317, 8'd205}: color_data = 12'h330;
			{9'd317, 8'd206}: color_data = 12'h9b0;
			{9'd317, 8'd207}: color_data = 12'hbc3;
			{9'd317, 8'd208}: color_data = 12'hffe;
			{9'd317, 8'd209}: color_data = 12'hffd;
			{9'd317, 8'd210}: color_data = 12'hac2;
			{9'd317, 8'd211}: color_data = 12'h9b0;
			{9'd317, 8'd212}: color_data = 12'h9b0;
			{9'd317, 8'd213}: color_data = 12'h9b0;
			{9'd317, 8'd214}: color_data = 12'h780;
			{9'd317, 8'd215}: color_data = 12'h230;
			{9'd317, 8'd216}: color_data = 12'h030;
			{9'd317, 8'd217}: color_data = 12'h140;
			{9'd317, 8'd218}: color_data = 12'h450;
			{9'd317, 8'd219}: color_data = 12'h770;
			{9'd317, 8'd220}: color_data = 12'h440;
			{9'd317, 8'd221}: color_data = 12'h000;
			{9'd317, 8'd222}: color_data = 12'h410;
			{9'd317, 8'd223}: color_data = 12'hd30;
			{9'd317, 8'd224}: color_data = 12'ha00;
			{9'd317, 8'd225}: color_data = 12'h700;
			{9'd317, 8'd226}: color_data = 12'h200;
			{9'd317, 8'd227}: color_data = 12'h700;
			{9'd317, 8'd228}: color_data = 12'hb00;
			{9'd317, 8'd229}: color_data = 12'ha00;
			{9'd317, 8'd230}: color_data = 12'h300;
			{9'd317, 8'd231}: color_data = 12'h820;
			{9'd317, 8'd232}: color_data = 12'hd20;
			{9'd317, 8'd233}: color_data = 12'h900;
			{9'd317, 8'd234}: color_data = 12'h500;
			{9'd317, 8'd235}: color_data = 12'h300;
			{9'd317, 8'd236}: color_data = 12'h900;
			{9'd317, 8'd237}: color_data = 12'hb00;
			{9'd317, 8'd238}: color_data = 12'h800;
			{9'd317, 8'd239}: color_data = 12'h100;
			{9'd318, 8'd24}: color_data = 12'h000;
			{9'd318, 8'd25}: color_data = 12'h000;
			{9'd318, 8'd26}: color_data = 12'h000;
			{9'd318, 8'd27}: color_data = 12'h000;
			{9'd318, 8'd28}: color_data = 12'h000;
			{9'd318, 8'd29}: color_data = 12'h000;
			{9'd318, 8'd30}: color_data = 12'h000;
			{9'd318, 8'd31}: color_data = 12'h000;
			{9'd318, 8'd32}: color_data = 12'h000;
			{9'd318, 8'd33}: color_data = 12'h000;
			{9'd318, 8'd34}: color_data = 12'h000;
			{9'd318, 8'd35}: color_data = 12'h000;
			{9'd318, 8'd36}: color_data = 12'h000;
			{9'd318, 8'd37}: color_data = 12'h000;
			{9'd318, 8'd38}: color_data = 12'h000;
			{9'd318, 8'd39}: color_data = 12'h000;
			{9'd318, 8'd40}: color_data = 12'h000;
			{9'd318, 8'd41}: color_data = 12'h000;
			{9'd318, 8'd42}: color_data = 12'h000;
			{9'd318, 8'd43}: color_data = 12'h000;
			{9'd318, 8'd45}: color_data = 12'h111;
			{9'd318, 8'd46}: color_data = 12'h888;
			{9'd318, 8'd47}: color_data = 12'h783;
			{9'd318, 8'd48}: color_data = 12'h670;
			{9'd318, 8'd49}: color_data = 12'h670;
			{9'd318, 8'd50}: color_data = 12'h220;
			{9'd318, 8'd51}: color_data = 12'h450;
			{9'd318, 8'd52}: color_data = 12'h9b0;
			{9'd318, 8'd53}: color_data = 12'hcd7;
			{9'd318, 8'd54}: color_data = 12'hfff;
			{9'd318, 8'd55}: color_data = 12'hdea;
			{9'd318, 8'd56}: color_data = 12'h9b0;
			{9'd318, 8'd57}: color_data = 12'h9b0;
			{9'd318, 8'd58}: color_data = 12'h9a0;
			{9'd318, 8'd59}: color_data = 12'h560;
			{9'd318, 8'd60}: color_data = 12'h020;
			{9'd318, 8'd61}: color_data = 12'h130;
			{9'd318, 8'd62}: color_data = 12'h240;
			{9'd318, 8'd63}: color_data = 12'h560;
			{9'd318, 8'd64}: color_data = 12'h760;
			{9'd318, 8'd65}: color_data = 12'h220;
			{9'd318, 8'd68}: color_data = 12'h036;
			{9'd318, 8'd69}: color_data = 12'h058;
			{9'd318, 8'd70}: color_data = 12'h002;
			{9'd318, 8'd71}: color_data = 12'h005;
			{9'd318, 8'd72}: color_data = 12'h005;
			{9'd318, 8'd73}: color_data = 12'h005;
			{9'd318, 8'd74}: color_data = 12'h005;
			{9'd318, 8'd75}: color_data = 12'h016;
			{9'd318, 8'd76}: color_data = 12'h05a;
			{9'd318, 8'd77}: color_data = 12'h023;
			{9'd318, 8'd128}: color_data = 12'h036;
			{9'd318, 8'd129}: color_data = 12'h058;
			{9'd318, 8'd130}: color_data = 12'h002;
			{9'd318, 8'd131}: color_data = 12'h005;
			{9'd318, 8'd132}: color_data = 12'h005;
			{9'd318, 8'd133}: color_data = 12'h005;
			{9'd318, 8'd134}: color_data = 12'h005;
			{9'd318, 8'd135}: color_data = 12'h016;
			{9'd318, 8'd136}: color_data = 12'h05a;
			{9'd318, 8'd137}: color_data = 12'h023;
			{9'd318, 8'd170}: color_data = 12'h000;
			{9'd318, 8'd171}: color_data = 12'h047;
			{9'd318, 8'd172}: color_data = 12'h047;
			{9'd318, 8'd173}: color_data = 12'h002;
			{9'd318, 8'd174}: color_data = 12'h005;
			{9'd318, 8'd175}: color_data = 12'h005;
			{9'd318, 8'd176}: color_data = 12'h005;
			{9'd318, 8'd177}: color_data = 12'h004;
			{9'd318, 8'd178}: color_data = 12'h017;
			{9'd318, 8'd179}: color_data = 12'h05a;
			{9'd318, 8'd180}: color_data = 12'h012;
			{9'd318, 8'd205}: color_data = 12'h330;
			{9'd318, 8'd206}: color_data = 12'h9b0;
			{9'd318, 8'd207}: color_data = 12'hbc3;
			{9'd318, 8'd208}: color_data = 12'hffe;
			{9'd318, 8'd209}: color_data = 12'hffd;
			{9'd318, 8'd210}: color_data = 12'hac2;
			{9'd318, 8'd211}: color_data = 12'h9b0;
			{9'd318, 8'd212}: color_data = 12'h9b0;
			{9'd318, 8'd213}: color_data = 12'h9b0;
			{9'd318, 8'd214}: color_data = 12'h780;
			{9'd318, 8'd215}: color_data = 12'h230;
			{9'd318, 8'd216}: color_data = 12'h030;
			{9'd318, 8'd217}: color_data = 12'h140;
			{9'd318, 8'd218}: color_data = 12'h450;
			{9'd318, 8'd219}: color_data = 12'h770;
			{9'd318, 8'd220}: color_data = 12'h440;
			{9'd318, 8'd221}: color_data = 12'h000;
			{9'd318, 8'd222}: color_data = 12'h310;
			{9'd318, 8'd223}: color_data = 12'he30;
			{9'd318, 8'd224}: color_data = 12'hc10;
			{9'd318, 8'd225}: color_data = 12'h800;
			{9'd318, 8'd226}: color_data = 12'h200;
			{9'd318, 8'd227}: color_data = 12'h600;
			{9'd318, 8'd228}: color_data = 12'ha00;
			{9'd318, 8'd229}: color_data = 12'h900;
			{9'd318, 8'd230}: color_data = 12'h300;
			{9'd318, 8'd231}: color_data = 12'h820;
			{9'd318, 8'd232}: color_data = 12'he30;
			{9'd318, 8'd233}: color_data = 12'hb00;
			{9'd318, 8'd234}: color_data = 12'h500;
			{9'd318, 8'd235}: color_data = 12'h200;
			{9'd318, 8'd236}: color_data = 12'h900;
			{9'd318, 8'd237}: color_data = 12'ha00;
			{9'd318, 8'd238}: color_data = 12'h700;
			{9'd318, 8'd239}: color_data = 12'h100;
			{9'd319, 8'd45}: color_data = 12'h000;
			{9'd319, 8'd46}: color_data = 12'h000;
			{9'd319, 8'd47}: color_data = 12'h000;
			{9'd319, 8'd48}: color_data = 12'h000;
			{9'd319, 8'd49}: color_data = 12'h000;
			{9'd319, 8'd50}: color_data = 12'h000;
			{9'd319, 8'd51}: color_data = 12'h560;
			{9'd319, 8'd52}: color_data = 12'h9b0;
			{9'd319, 8'd53}: color_data = 12'hcd7;
			{9'd319, 8'd54}: color_data = 12'hfff;
			{9'd319, 8'd55}: color_data = 12'hdea;
			{9'd319, 8'd56}: color_data = 12'h9b0;
			{9'd319, 8'd57}: color_data = 12'h9b0;
			{9'd319, 8'd58}: color_data = 12'h9a0;
			{9'd319, 8'd59}: color_data = 12'h560;
			{9'd319, 8'd60}: color_data = 12'h020;
			{9'd319, 8'd61}: color_data = 12'h130;
			{9'd319, 8'd62}: color_data = 12'h240;
			{9'd319, 8'd63}: color_data = 12'h560;
			{9'd319, 8'd64}: color_data = 12'h760;
			{9'd319, 8'd65}: color_data = 12'h220;
			{9'd319, 8'd68}: color_data = 12'h002;
			{9'd319, 8'd69}: color_data = 12'h005;
			{9'd319, 8'd70}: color_data = 12'h005;
			{9'd319, 8'd71}: color_data = 12'h005;
			{9'd319, 8'd72}: color_data = 12'h005;
			{9'd319, 8'd73}: color_data = 12'h005;
			{9'd319, 8'd74}: color_data = 12'h005;
			{9'd319, 8'd75}: color_data = 12'h005;
			{9'd319, 8'd76}: color_data = 12'h005;
			{9'd319, 8'd77}: color_data = 12'h001;
			{9'd319, 8'd128}: color_data = 12'h002;
			{9'd319, 8'd129}: color_data = 12'h005;
			{9'd319, 8'd130}: color_data = 12'h005;
			{9'd319, 8'd131}: color_data = 12'h005;
			{9'd319, 8'd132}: color_data = 12'h005;
			{9'd319, 8'd133}: color_data = 12'h005;
			{9'd319, 8'd134}: color_data = 12'h005;
			{9'd319, 8'd135}: color_data = 12'h005;
			{9'd319, 8'd136}: color_data = 12'h005;
			{9'd319, 8'd137}: color_data = 12'h001;
			{9'd319, 8'd170}: color_data = 12'h000;
			{9'd319, 8'd171}: color_data = 12'h003;
			{9'd319, 8'd172}: color_data = 12'h005;
			{9'd319, 8'd173}: color_data = 12'h005;
			{9'd319, 8'd174}: color_data = 12'h005;
			{9'd319, 8'd175}: color_data = 12'h005;
			{9'd319, 8'd176}: color_data = 12'h005;
			{9'd319, 8'd177}: color_data = 12'h005;
			{9'd319, 8'd178}: color_data = 12'h005;
			{9'd319, 8'd179}: color_data = 12'h004;
			{9'd319, 8'd180}: color_data = 12'h000;
			{9'd319, 8'd205}: color_data = 12'h330;
			{9'd319, 8'd206}: color_data = 12'h9b0;
			{9'd319, 8'd207}: color_data = 12'hbc3;
			{9'd319, 8'd208}: color_data = 12'hffe;
			{9'd319, 8'd209}: color_data = 12'hffd;
			{9'd319, 8'd210}: color_data = 12'hac2;
			{9'd319, 8'd211}: color_data = 12'h9b0;
			{9'd319, 8'd212}: color_data = 12'h9b0;
			{9'd319, 8'd213}: color_data = 12'h9b0;
			{9'd319, 8'd214}: color_data = 12'h780;
			{9'd319, 8'd215}: color_data = 12'h230;
			{9'd319, 8'd216}: color_data = 12'h030;
			{9'd319, 8'd217}: color_data = 12'h140;
			{9'd319, 8'd218}: color_data = 12'h450;
			{9'd319, 8'd219}: color_data = 12'h770;
			{9'd319, 8'd220}: color_data = 12'h440;
			{9'd319, 8'd221}: color_data = 12'h000;
			{9'd319, 8'd222}: color_data = 12'h300;
			{9'd319, 8'd223}: color_data = 12'he40;
			{9'd319, 8'd224}: color_data = 12'hf40;
			{9'd319, 8'd225}: color_data = 12'h800;
			{9'd319, 8'd226}: color_data = 12'h100;
			{9'd319, 8'd227}: color_data = 12'h600;
			{9'd319, 8'd228}: color_data = 12'ha00;
			{9'd319, 8'd229}: color_data = 12'h900;
			{9'd319, 8'd230}: color_data = 12'h300;
			{9'd319, 8'd231}: color_data = 12'h820;
			{9'd319, 8'd232}: color_data = 12'hf40;
			{9'd319, 8'd233}: color_data = 12'hd20;
			{9'd319, 8'd234}: color_data = 12'h400;
			{9'd319, 8'd235}: color_data = 12'h200;
			{9'd319, 8'd236}: color_data = 12'h900;
			{9'd319, 8'd237}: color_data = 12'ha00;
			{9'd319, 8'd238}: color_data = 12'h700;
			{9'd319, 8'd239}: color_data = 12'h100;
            default: color_data = 12'h3b9;
        endcase
endmodule
