module ending_rom(
        input wire clk,
        input wire [7:0] x,
        input wire [7:0] y,
        output reg [11:0] color_data
);

    (* rom_style = "block" *)

    //signal declaration
    reg [7:0] x_reg;
    reg [7:0] y_reg;

    always @(posedge clk) begin
        x_reg <= x;
        y_reg <= y;
    end

    always @*
        case ({x_reg, y_reg})
			// right: 8'd139, bottom: 8'd159
			{8'd1, 8'd26}: color_data = 12'hfc5;
			{8'd1, 8'd27}: color_data = 12'heb4;
			{8'd2, 8'd25}: color_data = 12'hfc4;
			{8'd2, 8'd26}: color_data = 12'hfc4;
			{8'd2, 8'd27}: color_data = 12'hfc4;
			{8'd2, 8'd28}: color_data = 12'hfc5;
			{8'd2, 8'd29}: color_data = 12'hfc5;
			{8'd2, 8'd30}: color_data = 12'hdb3;
			{8'd3, 8'd24}: color_data = 12'hfc5;
			{8'd3, 8'd25}: color_data = 12'hfc5;
			{8'd3, 8'd26}: color_data = 12'hfc5;
			{8'd3, 8'd27}: color_data = 12'hfc5;
			{8'd3, 8'd28}: color_data = 12'hfc5;
			{8'd3, 8'd29}: color_data = 12'hfc5;
			{8'd3, 8'd30}: color_data = 12'hfc5;
			{8'd3, 8'd31}: color_data = 12'hfc4;
			{8'd3, 8'd32}: color_data = 12'hfc4;
			{8'd3, 8'd33}: color_data = 12'hfb3;
			{8'd4, 8'd24}: color_data = 12'hfc5;
			{8'd4, 8'd25}: color_data = 12'hfc5;
			{8'd4, 8'd26}: color_data = 12'hfb3;
			{8'd4, 8'd27}: color_data = 12'hea1;
			{8'd4, 8'd28}: color_data = 12'heb2;
			{8'd4, 8'd29}: color_data = 12'hfc4;
			{8'd4, 8'd30}: color_data = 12'hfc5;
			{8'd4, 8'd31}: color_data = 12'hfc5;
			{8'd4, 8'd32}: color_data = 12'hfc4;
			{8'd4, 8'd33}: color_data = 12'hfc4;
			{8'd4, 8'd34}: color_data = 12'hfc5;
			{8'd4, 8'd35}: color_data = 12'hfc5;
			{8'd4, 8'd36}: color_data = 12'hdb3;
			{8'd5, 8'd23}: color_data = 12'hfd7;
			{8'd5, 8'd24}: color_data = 12'hfc5;
			{8'd5, 8'd25}: color_data = 12'hfc5;
			{8'd5, 8'd26}: color_data = 12'hea1;
			{8'd5, 8'd27}: color_data = 12'hd90;
			{8'd5, 8'd28}: color_data = 12'hd90;
			{8'd5, 8'd29}: color_data = 12'hd90;
			{8'd5, 8'd30}: color_data = 12'hea1;
			{8'd5, 8'd31}: color_data = 12'heb2;
			{8'd5, 8'd32}: color_data = 12'hfc4;
			{8'd5, 8'd33}: color_data = 12'hfc5;
			{8'd5, 8'd34}: color_data = 12'hfc5;
			{8'd5, 8'd35}: color_data = 12'hfc5;
			{8'd5, 8'd36}: color_data = 12'hfc5;
			{8'd5, 8'd37}: color_data = 12'hfc5;
			{8'd5, 8'd38}: color_data = 12'hec5;
			{8'd5, 8'd39}: color_data = 12'hfb3;
			{8'd6, 8'd23}: color_data = 12'hfc5;
			{8'd6, 8'd24}: color_data = 12'hfc5;
			{8'd6, 8'd25}: color_data = 12'hfc3;
			{8'd6, 8'd26}: color_data = 12'hd90;
			{8'd6, 8'd27}: color_data = 12'hd90;
			{8'd6, 8'd28}: color_data = 12'hd90;
			{8'd6, 8'd29}: color_data = 12'hd90;
			{8'd6, 8'd30}: color_data = 12'hd90;
			{8'd6, 8'd31}: color_data = 12'hd90;
			{8'd6, 8'd32}: color_data = 12'hd90;
			{8'd6, 8'd33}: color_data = 12'hea1;
			{8'd6, 8'd34}: color_data = 12'heb3;
			{8'd6, 8'd35}: color_data = 12'hfc4;
			{8'd6, 8'd36}: color_data = 12'hfc5;
			{8'd6, 8'd37}: color_data = 12'hfc5;
			{8'd6, 8'd38}: color_data = 12'hfc5;
			{8'd6, 8'd39}: color_data = 12'hfc5;
			{8'd6, 8'd40}: color_data = 12'hfc4;
			{8'd6, 8'd77}: color_data = 12'h000;
			{8'd6, 8'd78}: color_data = 12'h000;
			{8'd6, 8'd79}: color_data = 12'h000;
			{8'd6, 8'd80}: color_data = 12'h000;
			{8'd7, 8'd23}: color_data = 12'hfc4;
			{8'd7, 8'd24}: color_data = 12'hfc5;
			{8'd7, 8'd25}: color_data = 12'hea2;
			{8'd7, 8'd26}: color_data = 12'hd90;
			{8'd7, 8'd27}: color_data = 12'hd90;
			{8'd7, 8'd28}: color_data = 12'hd90;
			{8'd7, 8'd29}: color_data = 12'hd90;
			{8'd7, 8'd30}: color_data = 12'hd90;
			{8'd7, 8'd31}: color_data = 12'hd90;
			{8'd7, 8'd32}: color_data = 12'hd90;
			{8'd7, 8'd33}: color_data = 12'hd90;
			{8'd7, 8'd34}: color_data = 12'hd90;
			{8'd7, 8'd35}: color_data = 12'hd90;
			{8'd7, 8'd36}: color_data = 12'hea1;
			{8'd7, 8'd37}: color_data = 12'heb2;
			{8'd7, 8'd38}: color_data = 12'hfc4;
			{8'd7, 8'd39}: color_data = 12'hfc5;
			{8'd7, 8'd40}: color_data = 12'hfc5;
			{8'd7, 8'd41}: color_data = 12'hfc6;
			{8'd7, 8'd75}: color_data = 12'h000;
			{8'd7, 8'd76}: color_data = 12'h020;
			{8'd7, 8'd77}: color_data = 12'h062;
			{8'd7, 8'd78}: color_data = 12'h082;
			{8'd7, 8'd79}: color_data = 12'h072;
			{8'd7, 8'd80}: color_data = 12'h041;
			{8'd7, 8'd81}: color_data = 12'h000;
			{8'd8, 8'd22}: color_data = 12'hfd6;
			{8'd8, 8'd23}: color_data = 12'hfc5;
			{8'd8, 8'd24}: color_data = 12'hfc4;
			{8'd8, 8'd25}: color_data = 12'heb3;
			{8'd8, 8'd26}: color_data = 12'hea1;
			{8'd8, 8'd27}: color_data = 12'hda0;
			{8'd8, 8'd28}: color_data = 12'hd90;
			{8'd8, 8'd29}: color_data = 12'hd90;
			{8'd8, 8'd30}: color_data = 12'hd90;
			{8'd8, 8'd31}: color_data = 12'hd90;
			{8'd8, 8'd32}: color_data = 12'hd90;
			{8'd8, 8'd33}: color_data = 12'hd90;
			{8'd8, 8'd34}: color_data = 12'hd90;
			{8'd8, 8'd35}: color_data = 12'hd90;
			{8'd8, 8'd36}: color_data = 12'hd90;
			{8'd8, 8'd37}: color_data = 12'hd90;
			{8'd8, 8'd38}: color_data = 12'hea0;
			{8'd8, 8'd39}: color_data = 12'hfc5;
			{8'd8, 8'd40}: color_data = 12'hfc5;
			{8'd8, 8'd41}: color_data = 12'hfc6;
			{8'd8, 8'd74}: color_data = 12'h000;
			{8'd8, 8'd75}: color_data = 12'h031;
			{8'd8, 8'd76}: color_data = 12'h093;
			{8'd8, 8'd77}: color_data = 12'h0a4;
			{8'd8, 8'd78}: color_data = 12'h0a3;
			{8'd8, 8'd79}: color_data = 12'h0a3;
			{8'd8, 8'd80}: color_data = 12'h0a3;
			{8'd8, 8'd81}: color_data = 12'h041;
			{8'd8, 8'd82}: color_data = 12'h000;
			{8'd9, 8'd23}: color_data = 12'hfc5;
			{8'd9, 8'd24}: color_data = 12'hfc5;
			{8'd9, 8'd25}: color_data = 12'hfc5;
			{8'd9, 8'd26}: color_data = 12'hfc5;
			{8'd9, 8'd27}: color_data = 12'hfc4;
			{8'd9, 8'd28}: color_data = 12'hfb4;
			{8'd9, 8'd29}: color_data = 12'hfb3;
			{8'd9, 8'd30}: color_data = 12'hea0;
			{8'd9, 8'd31}: color_data = 12'hd90;
			{8'd9, 8'd32}: color_data = 12'hd90;
			{8'd9, 8'd33}: color_data = 12'hd90;
			{8'd9, 8'd34}: color_data = 12'hd90;
			{8'd9, 8'd35}: color_data = 12'hd90;
			{8'd9, 8'd36}: color_data = 12'hd90;
			{8'd9, 8'd37}: color_data = 12'hd90;
			{8'd9, 8'd38}: color_data = 12'hda0;
			{8'd9, 8'd39}: color_data = 12'hfc4;
			{8'd9, 8'd40}: color_data = 12'hfc5;
			{8'd9, 8'd41}: color_data = 12'hec5;
			{8'd9, 8'd74}: color_data = 12'h031;
			{8'd9, 8'd75}: color_data = 12'h093;
			{8'd9, 8'd76}: color_data = 12'h0a3;
			{8'd9, 8'd77}: color_data = 12'h0a3;
			{8'd9, 8'd78}: color_data = 12'h0a3;
			{8'd9, 8'd79}: color_data = 12'h0a3;
			{8'd9, 8'd80}: color_data = 12'h0a3;
			{8'd9, 8'd81}: color_data = 12'h093;
			{8'd9, 8'd82}: color_data = 12'h020;
			{8'd10, 8'd22}: color_data = 12'hfd6;
			{8'd10, 8'd23}: color_data = 12'hfc5;
			{8'd10, 8'd24}: color_data = 12'hfc6;
			{8'd10, 8'd25}: color_data = 12'hfc6;
			{8'd10, 8'd26}: color_data = 12'hfc5;
			{8'd10, 8'd27}: color_data = 12'hfc5;
			{8'd10, 8'd28}: color_data = 12'hfc5;
			{8'd10, 8'd29}: color_data = 12'hfc6;
			{8'd10, 8'd30}: color_data = 12'hea1;
			{8'd10, 8'd31}: color_data = 12'hd90;
			{8'd10, 8'd32}: color_data = 12'hd90;
			{8'd10, 8'd33}: color_data = 12'hd90;
			{8'd10, 8'd34}: color_data = 12'hd90;
			{8'd10, 8'd35}: color_data = 12'hd90;
			{8'd10, 8'd36}: color_data = 12'hd90;
			{8'd10, 8'd37}: color_data = 12'hd90;
			{8'd10, 8'd38}: color_data = 12'hea1;
			{8'd10, 8'd39}: color_data = 12'hfc5;
			{8'd10, 8'd40}: color_data = 12'hfc4;
			{8'd10, 8'd73}: color_data = 12'h000;
			{8'd10, 8'd74}: color_data = 12'h072;
			{8'd10, 8'd75}: color_data = 12'h0a3;
			{8'd10, 8'd76}: color_data = 12'h0a3;
			{8'd10, 8'd77}: color_data = 12'h0a3;
			{8'd10, 8'd78}: color_data = 12'h0a3;
			{8'd10, 8'd79}: color_data = 12'h0a3;
			{8'd10, 8'd80}: color_data = 12'h0a3;
			{8'd10, 8'd81}: color_data = 12'h0a3;
			{8'd10, 8'd82}: color_data = 12'h041;
			{8'd11, 8'd22}: color_data = 12'hfc4;
			{8'd11, 8'd23}: color_data = 12'hfc4;
			{8'd11, 8'd24}: color_data = 12'hfc4;
			{8'd11, 8'd25}: color_data = 12'hfb3;
			{8'd11, 8'd26}: color_data = 12'hfc4;
			{8'd11, 8'd27}: color_data = 12'hfc5;
			{8'd11, 8'd28}: color_data = 12'hfc5;
			{8'd11, 8'd29}: color_data = 12'hfc4;
			{8'd11, 8'd30}: color_data = 12'hd90;
			{8'd11, 8'd31}: color_data = 12'hd90;
			{8'd11, 8'd32}: color_data = 12'hd90;
			{8'd11, 8'd33}: color_data = 12'hd90;
			{8'd11, 8'd34}: color_data = 12'heb2;
			{8'd11, 8'd35}: color_data = 12'hfb4;
			{8'd11, 8'd36}: color_data = 12'heb2;
			{8'd11, 8'd37}: color_data = 12'hea1;
			{8'd11, 8'd38}: color_data = 12'heb3;
			{8'd11, 8'd39}: color_data = 12'hfc5;
			{8'd11, 8'd40}: color_data = 12'hfc5;
			{8'd11, 8'd72}: color_data = 12'h000;
			{8'd11, 8'd73}: color_data = 12'h051;
			{8'd11, 8'd74}: color_data = 12'h0a3;
			{8'd11, 8'd75}: color_data = 12'h0a3;
			{8'd11, 8'd76}: color_data = 12'h0a3;
			{8'd11, 8'd77}: color_data = 12'h0a3;
			{8'd11, 8'd78}: color_data = 12'h0a3;
			{8'd11, 8'd79}: color_data = 12'h0a3;
			{8'd11, 8'd80}: color_data = 12'h0a3;
			{8'd11, 8'd81}: color_data = 12'h0a3;
			{8'd11, 8'd82}: color_data = 12'h041;
			{8'd11, 8'd102}: color_data = 12'h000;
			{8'd11, 8'd103}: color_data = 12'h000;
			{8'd11, 8'd104}: color_data = 12'h000;
			{8'd12, 8'd22}: color_data = 12'hfc4;
			{8'd12, 8'd23}: color_data = 12'hfc5;
			{8'd12, 8'd24}: color_data = 12'heb2;
			{8'd12, 8'd25}: color_data = 12'hd90;
			{8'd12, 8'd26}: color_data = 12'hd90;
			{8'd12, 8'd27}: color_data = 12'hda0;
			{8'd12, 8'd28}: color_data = 12'hea1;
			{8'd12, 8'd29}: color_data = 12'hea1;
			{8'd12, 8'd30}: color_data = 12'hd90;
			{8'd12, 8'd31}: color_data = 12'hd90;
			{8'd12, 8'd32}: color_data = 12'hd90;
			{8'd12, 8'd33}: color_data = 12'hea0;
			{8'd12, 8'd34}: color_data = 12'hfc5;
			{8'd12, 8'd35}: color_data = 12'hfc5;
			{8'd12, 8'd36}: color_data = 12'hfc5;
			{8'd12, 8'd37}: color_data = 12'hfc5;
			{8'd12, 8'd38}: color_data = 12'hfc5;
			{8'd12, 8'd39}: color_data = 12'hfc5;
			{8'd12, 8'd40}: color_data = 12'hfc5;
			{8'd12, 8'd72}: color_data = 12'h010;
			{8'd12, 8'd73}: color_data = 12'h083;
			{8'd12, 8'd74}: color_data = 12'h0a3;
			{8'd12, 8'd75}: color_data = 12'h0a3;
			{8'd12, 8'd76}: color_data = 12'h0a3;
			{8'd12, 8'd77}: color_data = 12'h0a3;
			{8'd12, 8'd78}: color_data = 12'h0a3;
			{8'd12, 8'd79}: color_data = 12'h0a3;
			{8'd12, 8'd80}: color_data = 12'h0a3;
			{8'd12, 8'd81}: color_data = 12'h0a3;
			{8'd12, 8'd82}: color_data = 12'h041;
			{8'd12, 8'd100}: color_data = 12'h000;
			{8'd12, 8'd101}: color_data = 12'h020;
			{8'd12, 8'd102}: color_data = 12'h062;
			{8'd12, 8'd103}: color_data = 12'h072;
			{8'd12, 8'd104}: color_data = 12'h062;
			{8'd12, 8'd105}: color_data = 12'h031;
			{8'd12, 8'd106}: color_data = 12'h000;
			{8'd13, 8'd22}: color_data = 12'hfc5;
			{8'd13, 8'd23}: color_data = 12'hfc5;
			{8'd13, 8'd24}: color_data = 12'hea1;
			{8'd13, 8'd25}: color_data = 12'hd90;
			{8'd13, 8'd26}: color_data = 12'hd90;
			{8'd13, 8'd27}: color_data = 12'hd90;
			{8'd13, 8'd28}: color_data = 12'hd90;
			{8'd13, 8'd29}: color_data = 12'hd90;
			{8'd13, 8'd30}: color_data = 12'hd90;
			{8'd13, 8'd31}: color_data = 12'hd90;
			{8'd13, 8'd32}: color_data = 12'hd90;
			{8'd13, 8'd33}: color_data = 12'hea0;
			{8'd13, 8'd34}: color_data = 12'hfc4;
			{8'd13, 8'd35}: color_data = 12'hfc5;
			{8'd13, 8'd36}: color_data = 12'hfc5;
			{8'd13, 8'd37}: color_data = 12'hfc5;
			{8'd13, 8'd38}: color_data = 12'hfc5;
			{8'd13, 8'd39}: color_data = 12'hfc5;
			{8'd13, 8'd40}: color_data = 12'hfd5;
			{8'd13, 8'd72}: color_data = 12'h051;
			{8'd13, 8'd73}: color_data = 12'h0a3;
			{8'd13, 8'd74}: color_data = 12'h0a3;
			{8'd13, 8'd75}: color_data = 12'h0a3;
			{8'd13, 8'd76}: color_data = 12'h0a3;
			{8'd13, 8'd77}: color_data = 12'h0a3;
			{8'd13, 8'd78}: color_data = 12'h0a3;
			{8'd13, 8'd79}: color_data = 12'h0a3;
			{8'd13, 8'd80}: color_data = 12'h0a3;
			{8'd13, 8'd81}: color_data = 12'h0a3;
			{8'd13, 8'd82}: color_data = 12'h041;
			{8'd13, 8'd99}: color_data = 12'h000;
			{8'd13, 8'd100}: color_data = 12'h041;
			{8'd13, 8'd101}: color_data = 12'h093;
			{8'd13, 8'd102}: color_data = 12'h0a4;
			{8'd13, 8'd103}: color_data = 12'h0a3;
			{8'd13, 8'd104}: color_data = 12'h0a4;
			{8'd13, 8'd105}: color_data = 12'h093;
			{8'd13, 8'd106}: color_data = 12'h031;
			{8'd14, 8'd22}: color_data = 12'hfc5;
			{8'd14, 8'd23}: color_data = 12'hfc5;
			{8'd14, 8'd24}: color_data = 12'hea0;
			{8'd14, 8'd25}: color_data = 12'hd90;
			{8'd14, 8'd26}: color_data = 12'hd90;
			{8'd14, 8'd27}: color_data = 12'hd90;
			{8'd14, 8'd28}: color_data = 12'hd90;
			{8'd14, 8'd29}: color_data = 12'hd90;
			{8'd14, 8'd30}: color_data = 12'hd90;
			{8'd14, 8'd31}: color_data = 12'hd90;
			{8'd14, 8'd32}: color_data = 12'hd90;
			{8'd14, 8'd33}: color_data = 12'hd90;
			{8'd14, 8'd34}: color_data = 12'hd90;
			{8'd14, 8'd35}: color_data = 12'hda0;
			{8'd14, 8'd36}: color_data = 12'hea1;
			{8'd14, 8'd37}: color_data = 12'hfb3;
			{8'd14, 8'd38}: color_data = 12'hfc5;
			{8'd14, 8'd39}: color_data = 12'hfc6;
			{8'd14, 8'd71}: color_data = 12'h000;
			{8'd14, 8'd72}: color_data = 12'h072;
			{8'd14, 8'd73}: color_data = 12'h0a3;
			{8'd14, 8'd74}: color_data = 12'h0a3;
			{8'd14, 8'd75}: color_data = 12'h0a3;
			{8'd14, 8'd76}: color_data = 12'h0a3;
			{8'd14, 8'd77}: color_data = 12'h0a3;
			{8'd14, 8'd78}: color_data = 12'h0a3;
			{8'd14, 8'd79}: color_data = 12'h0a3;
			{8'd14, 8'd80}: color_data = 12'h0a3;
			{8'd14, 8'd81}: color_data = 12'h093;
			{8'd14, 8'd82}: color_data = 12'h020;
			{8'd14, 8'd98}: color_data = 12'h000;
			{8'd14, 8'd99}: color_data = 12'h041;
			{8'd14, 8'd100}: color_data = 12'h0a3;
			{8'd14, 8'd101}: color_data = 12'h0a3;
			{8'd14, 8'd102}: color_data = 12'h0a3;
			{8'd14, 8'd103}: color_data = 12'h0a3;
			{8'd14, 8'd104}: color_data = 12'h0a3;
			{8'd14, 8'd105}: color_data = 12'h0a4;
			{8'd14, 8'd106}: color_data = 12'h072;
			{8'd14, 8'd107}: color_data = 12'h000;
			{8'd15, 8'd21}: color_data = 12'hec5;
			{8'd15, 8'd22}: color_data = 12'hfc5;
			{8'd15, 8'd23}: color_data = 12'hfc5;
			{8'd15, 8'd24}: color_data = 12'heb3;
			{8'd15, 8'd25}: color_data = 12'hea1;
			{8'd15, 8'd26}: color_data = 12'hda0;
			{8'd15, 8'd27}: color_data = 12'hd90;
			{8'd15, 8'd28}: color_data = 12'hd90;
			{8'd15, 8'd29}: color_data = 12'hd90;
			{8'd15, 8'd30}: color_data = 12'hd90;
			{8'd15, 8'd31}: color_data = 12'hd90;
			{8'd15, 8'd32}: color_data = 12'hd90;
			{8'd15, 8'd33}: color_data = 12'hd90;
			{8'd15, 8'd34}: color_data = 12'hd90;
			{8'd15, 8'd35}: color_data = 12'hd90;
			{8'd15, 8'd36}: color_data = 12'hd90;
			{8'd15, 8'd37}: color_data = 12'heb2;
			{8'd15, 8'd38}: color_data = 12'hfc5;
			{8'd15, 8'd39}: color_data = 12'hfc5;
			{8'd15, 8'd68}: color_data = 12'h000;
			{8'd15, 8'd69}: color_data = 12'h000;
			{8'd15, 8'd70}: color_data = 12'h000;
			{8'd15, 8'd71}: color_data = 12'h010;
			{8'd15, 8'd72}: color_data = 12'h052;
			{8'd15, 8'd73}: color_data = 12'h093;
			{8'd15, 8'd74}: color_data = 12'h0a3;
			{8'd15, 8'd75}: color_data = 12'h0a3;
			{8'd15, 8'd76}: color_data = 12'h0a3;
			{8'd15, 8'd77}: color_data = 12'h0a3;
			{8'd15, 8'd78}: color_data = 12'h0a3;
			{8'd15, 8'd79}: color_data = 12'h0a3;
			{8'd15, 8'd80}: color_data = 12'h0a4;
			{8'd15, 8'd81}: color_data = 12'h062;
			{8'd15, 8'd82}: color_data = 12'h000;
			{8'd15, 8'd98}: color_data = 12'h010;
			{8'd15, 8'd99}: color_data = 12'h083;
			{8'd15, 8'd100}: color_data = 12'h0a3;
			{8'd15, 8'd101}: color_data = 12'h0a3;
			{8'd15, 8'd102}: color_data = 12'h0a3;
			{8'd15, 8'd103}: color_data = 12'h0a3;
			{8'd15, 8'd104}: color_data = 12'h0a3;
			{8'd15, 8'd105}: color_data = 12'h0a3;
			{8'd15, 8'd106}: color_data = 12'h083;
			{8'd15, 8'd107}: color_data = 12'h000;
			{8'd15, 8'd140}: color_data = 12'h000;
			{8'd15, 8'd141}: color_data = 12'h100;
			{8'd15, 8'd142}: color_data = 12'h211;
			{8'd15, 8'd143}: color_data = 12'h100;
			{8'd15, 8'd144}: color_data = 12'h111;
			{8'd15, 8'd145}: color_data = 12'h000;
			{8'd16, 8'd21}: color_data = 12'hfc5;
			{8'd16, 8'd22}: color_data = 12'hfc5;
			{8'd16, 8'd23}: color_data = 12'hfc6;
			{8'd16, 8'd24}: color_data = 12'hfc6;
			{8'd16, 8'd25}: color_data = 12'hfc6;
			{8'd16, 8'd26}: color_data = 12'hfc5;
			{8'd16, 8'd27}: color_data = 12'hfc4;
			{8'd16, 8'd28}: color_data = 12'heb2;
			{8'd16, 8'd29}: color_data = 12'hea1;
			{8'd16, 8'd30}: color_data = 12'hd90;
			{8'd16, 8'd31}: color_data = 12'hd90;
			{8'd16, 8'd32}: color_data = 12'hd90;
			{8'd16, 8'd33}: color_data = 12'hd90;
			{8'd16, 8'd34}: color_data = 12'hd90;
			{8'd16, 8'd35}: color_data = 12'hd90;
			{8'd16, 8'd36}: color_data = 12'hd90;
			{8'd16, 8'd37}: color_data = 12'hfb3;
			{8'd16, 8'd38}: color_data = 12'hfc5;
			{8'd16, 8'd39}: color_data = 12'hfc4;
			{8'd16, 8'd63}: color_data = 12'h000;
			{8'd16, 8'd64}: color_data = 12'h000;
			{8'd16, 8'd65}: color_data = 12'h020;
			{8'd16, 8'd66}: color_data = 12'h041;
			{8'd16, 8'd67}: color_data = 12'h051;
			{8'd16, 8'd68}: color_data = 12'h062;
			{8'd16, 8'd69}: color_data = 12'h072;
			{8'd16, 8'd70}: color_data = 12'h083;
			{8'd16, 8'd71}: color_data = 12'h083;
			{8'd16, 8'd72}: color_data = 12'h072;
			{8'd16, 8'd73}: color_data = 12'h0a3;
			{8'd16, 8'd74}: color_data = 12'h0a3;
			{8'd16, 8'd75}: color_data = 12'h0a3;
			{8'd16, 8'd76}: color_data = 12'h0a3;
			{8'd16, 8'd77}: color_data = 12'h0a3;
			{8'd16, 8'd78}: color_data = 12'h0a3;
			{8'd16, 8'd79}: color_data = 12'h0a3;
			{8'd16, 8'd80}: color_data = 12'h082;
			{8'd16, 8'd81}: color_data = 12'h010;
			{8'd16, 8'd98}: color_data = 12'h041;
			{8'd16, 8'd99}: color_data = 12'h0a3;
			{8'd16, 8'd100}: color_data = 12'h0a3;
			{8'd16, 8'd101}: color_data = 12'h0a3;
			{8'd16, 8'd102}: color_data = 12'h0a3;
			{8'd16, 8'd103}: color_data = 12'h0a3;
			{8'd16, 8'd104}: color_data = 12'h0a3;
			{8'd16, 8'd105}: color_data = 12'h0a3;
			{8'd16, 8'd106}: color_data = 12'h072;
			{8'd16, 8'd107}: color_data = 12'h000;
			{8'd16, 8'd139}: color_data = 12'h000;
			{8'd16, 8'd140}: color_data = 12'h321;
			{8'd16, 8'd141}: color_data = 12'h533;
			{8'd16, 8'd142}: color_data = 12'h643;
			{8'd16, 8'd143}: color_data = 12'h532;
			{8'd16, 8'd144}: color_data = 12'h643;
			{8'd16, 8'd145}: color_data = 12'h653;
			{8'd16, 8'd146}: color_data = 12'h000;
			{8'd17, 8'd20}: color_data = 12'hfc5;
			{8'd17, 8'd21}: color_data = 12'hfc4;
			{8'd17, 8'd22}: color_data = 12'hfc5;
			{8'd17, 8'd23}: color_data = 12'hfb2;
			{8'd17, 8'd24}: color_data = 12'heb2;
			{8'd17, 8'd25}: color_data = 12'heb2;
			{8'd17, 8'd26}: color_data = 12'heb2;
			{8'd17, 8'd27}: color_data = 12'heb2;
			{8'd17, 8'd28}: color_data = 12'heb3;
			{8'd17, 8'd29}: color_data = 12'hfc4;
			{8'd17, 8'd30}: color_data = 12'hfc4;
			{8'd17, 8'd31}: color_data = 12'hfb3;
			{8'd17, 8'd32}: color_data = 12'heb2;
			{8'd17, 8'd33}: color_data = 12'hea1;
			{8'd17, 8'd34}: color_data = 12'hd90;
			{8'd17, 8'd35}: color_data = 12'hd90;
			{8'd17, 8'd36}: color_data = 12'hd90;
			{8'd17, 8'd37}: color_data = 12'hfb3;
			{8'd17, 8'd38}: color_data = 12'hfc5;
			{8'd17, 8'd39}: color_data = 12'hfc4;
			{8'd17, 8'd61}: color_data = 12'h000;
			{8'd17, 8'd62}: color_data = 12'h031;
			{8'd17, 8'd63}: color_data = 12'h062;
			{8'd17, 8'd64}: color_data = 12'h083;
			{8'd17, 8'd65}: color_data = 12'h093;
			{8'd17, 8'd66}: color_data = 12'h0a3;
			{8'd17, 8'd67}: color_data = 12'h0a3;
			{8'd17, 8'd68}: color_data = 12'h0a3;
			{8'd17, 8'd69}: color_data = 12'h0a3;
			{8'd17, 8'd70}: color_data = 12'h0a3;
			{8'd17, 8'd71}: color_data = 12'h0a3;
			{8'd17, 8'd72}: color_data = 12'h0a3;
			{8'd17, 8'd73}: color_data = 12'h0a3;
			{8'd17, 8'd74}: color_data = 12'h0a3;
			{8'd17, 8'd75}: color_data = 12'h0a3;
			{8'd17, 8'd76}: color_data = 12'h0a3;
			{8'd17, 8'd77}: color_data = 12'h0a3;
			{8'd17, 8'd78}: color_data = 12'h0a3;
			{8'd17, 8'd79}: color_data = 12'h093;
			{8'd17, 8'd80}: color_data = 12'h431;
			{8'd17, 8'd81}: color_data = 12'h310;
			{8'd17, 8'd82}: color_data = 12'h000;
			{8'd17, 8'd83}: color_data = 12'h000;
			{8'd17, 8'd84}: color_data = 12'h000;
			{8'd17, 8'd97}: color_data = 12'h000;
			{8'd17, 8'd98}: color_data = 12'h062;
			{8'd17, 8'd99}: color_data = 12'h0a4;
			{8'd17, 8'd100}: color_data = 12'h0a3;
			{8'd17, 8'd101}: color_data = 12'h0a3;
			{8'd17, 8'd102}: color_data = 12'h0a3;
			{8'd17, 8'd103}: color_data = 12'h0a3;
			{8'd17, 8'd104}: color_data = 12'h0a3;
			{8'd17, 8'd105}: color_data = 12'h0a3;
			{8'd17, 8'd106}: color_data = 12'h051;
			{8'd17, 8'd138}: color_data = 12'h100;
			{8'd17, 8'd139}: color_data = 12'h422;
			{8'd17, 8'd140}: color_data = 12'h643;
			{8'd17, 8'd141}: color_data = 12'h643;
			{8'd17, 8'd142}: color_data = 12'h633;
			{8'd17, 8'd143}: color_data = 12'h643;
			{8'd17, 8'd144}: color_data = 12'h532;
			{8'd17, 8'd145}: color_data = 12'h974;
			{8'd17, 8'd146}: color_data = 12'h000;
			{8'd18, 8'd20}: color_data = 12'hfc6;
			{8'd18, 8'd21}: color_data = 12'hfc5;
			{8'd18, 8'd22}: color_data = 12'hfc4;
			{8'd18, 8'd23}: color_data = 12'hd90;
			{8'd18, 8'd24}: color_data = 12'hd90;
			{8'd18, 8'd25}: color_data = 12'hd90;
			{8'd18, 8'd26}: color_data = 12'hd90;
			{8'd18, 8'd27}: color_data = 12'hd90;
			{8'd18, 8'd28}: color_data = 12'hd90;
			{8'd18, 8'd29}: color_data = 12'hd90;
			{8'd18, 8'd30}: color_data = 12'hea1;
			{8'd18, 8'd31}: color_data = 12'heb2;
			{8'd18, 8'd32}: color_data = 12'hfc5;
			{8'd18, 8'd33}: color_data = 12'hfc5;
			{8'd18, 8'd34}: color_data = 12'hfc5;
			{8'd18, 8'd35}: color_data = 12'hfb4;
			{8'd18, 8'd36}: color_data = 12'heb2;
			{8'd18, 8'd37}: color_data = 12'hfc5;
			{8'd18, 8'd38}: color_data = 12'hfc5;
			{8'd18, 8'd39}: color_data = 12'hfc5;
			{8'd18, 8'd59}: color_data = 12'h000;
			{8'd18, 8'd60}: color_data = 12'h031;
			{8'd18, 8'd61}: color_data = 12'h072;
			{8'd18, 8'd62}: color_data = 12'h0a3;
			{8'd18, 8'd63}: color_data = 12'h0a4;
			{8'd18, 8'd64}: color_data = 12'h0a3;
			{8'd18, 8'd65}: color_data = 12'h0a3;
			{8'd18, 8'd66}: color_data = 12'h0a3;
			{8'd18, 8'd67}: color_data = 12'h0a3;
			{8'd18, 8'd68}: color_data = 12'h0a3;
			{8'd18, 8'd69}: color_data = 12'h0a3;
			{8'd18, 8'd70}: color_data = 12'h0a3;
			{8'd18, 8'd71}: color_data = 12'h0a3;
			{8'd18, 8'd72}: color_data = 12'h0a3;
			{8'd18, 8'd73}: color_data = 12'h0a3;
			{8'd18, 8'd74}: color_data = 12'h0a3;
			{8'd18, 8'd75}: color_data = 12'h0a3;
			{8'd18, 8'd76}: color_data = 12'h0a3;
			{8'd18, 8'd77}: color_data = 12'h0a3;
			{8'd18, 8'd78}: color_data = 12'h093;
			{8'd18, 8'd79}: color_data = 12'h331;
			{8'd18, 8'd80}: color_data = 12'h632;
			{8'd18, 8'd81}: color_data = 12'h876;
			{8'd18, 8'd82}: color_data = 12'hca8;
			{8'd18, 8'd83}: color_data = 12'hca9;
			{8'd18, 8'd84}: color_data = 12'ha87;
			{8'd18, 8'd85}: color_data = 12'h543;
			{8'd18, 8'd86}: color_data = 12'h000;
			{8'd18, 8'd97}: color_data = 12'h000;
			{8'd18, 8'd98}: color_data = 12'h072;
			{8'd18, 8'd99}: color_data = 12'h0b4;
			{8'd18, 8'd100}: color_data = 12'h0a3;
			{8'd18, 8'd101}: color_data = 12'h093;
			{8'd18, 8'd102}: color_data = 12'h083;
			{8'd18, 8'd103}: color_data = 12'h174;
			{8'd18, 8'd104}: color_data = 12'h385;
			{8'd18, 8'd105}: color_data = 12'h374;
			{8'd18, 8'd106}: color_data = 12'h132;
			{8'd18, 8'd107}: color_data = 12'h000;
			{8'd18, 8'd130}: color_data = 12'h000;
			{8'd18, 8'd131}: color_data = 12'h000;
			{8'd18, 8'd132}: color_data = 12'h001;
			{8'd18, 8'd133}: color_data = 12'h001;
			{8'd18, 8'd134}: color_data = 12'h000;
			{8'd18, 8'd137}: color_data = 12'h000;
			{8'd18, 8'd138}: color_data = 12'h322;
			{8'd18, 8'd139}: color_data = 12'h643;
			{8'd18, 8'd140}: color_data = 12'h633;
			{8'd18, 8'd141}: color_data = 12'h633;
			{8'd18, 8'd142}: color_data = 12'h633;
			{8'd18, 8'd143}: color_data = 12'h643;
			{8'd18, 8'd144}: color_data = 12'h532;
			{8'd18, 8'd145}: color_data = 12'h763;
			{8'd18, 8'd146}: color_data = 12'h432;
			{8'd19, 8'd20}: color_data = 12'hfc5;
			{8'd19, 8'd21}: color_data = 12'hfc5;
			{8'd19, 8'd22}: color_data = 12'hfb3;
			{8'd19, 8'd23}: color_data = 12'hd90;
			{8'd19, 8'd24}: color_data = 12'hd90;
			{8'd19, 8'd25}: color_data = 12'hd90;
			{8'd19, 8'd26}: color_data = 12'hd90;
			{8'd19, 8'd27}: color_data = 12'hd90;
			{8'd19, 8'd28}: color_data = 12'hd90;
			{8'd19, 8'd29}: color_data = 12'hd90;
			{8'd19, 8'd30}: color_data = 12'hd90;
			{8'd19, 8'd31}: color_data = 12'hd90;
			{8'd19, 8'd32}: color_data = 12'hd90;
			{8'd19, 8'd33}: color_data = 12'hda0;
			{8'd19, 8'd34}: color_data = 12'heb2;
			{8'd19, 8'd35}: color_data = 12'hfc5;
			{8'd19, 8'd36}: color_data = 12'hfc5;
			{8'd19, 8'd37}: color_data = 12'hfc5;
			{8'd19, 8'd38}: color_data = 12'hfc4;
			{8'd19, 8'd39}: color_data = 12'hfff;
			{8'd19, 8'd57}: color_data = 12'h000;
			{8'd19, 8'd58}: color_data = 12'h010;
			{8'd19, 8'd59}: color_data = 12'h062;
			{8'd19, 8'd60}: color_data = 12'h0a3;
			{8'd19, 8'd61}: color_data = 12'h0a3;
			{8'd19, 8'd62}: color_data = 12'h0a3;
			{8'd19, 8'd63}: color_data = 12'h0a3;
			{8'd19, 8'd64}: color_data = 12'h0a3;
			{8'd19, 8'd65}: color_data = 12'h0a3;
			{8'd19, 8'd66}: color_data = 12'h0a3;
			{8'd19, 8'd67}: color_data = 12'h0a3;
			{8'd19, 8'd68}: color_data = 12'h0a3;
			{8'd19, 8'd69}: color_data = 12'h0a3;
			{8'd19, 8'd70}: color_data = 12'h0a3;
			{8'd19, 8'd71}: color_data = 12'h0a3;
			{8'd19, 8'd72}: color_data = 12'h0a3;
			{8'd19, 8'd73}: color_data = 12'h0a3;
			{8'd19, 8'd74}: color_data = 12'h0a3;
			{8'd19, 8'd75}: color_data = 12'h0a3;
			{8'd19, 8'd76}: color_data = 12'h0a3;
			{8'd19, 8'd77}: color_data = 12'h093;
			{8'd19, 8'd78}: color_data = 12'h241;
			{8'd19, 8'd79}: color_data = 12'h632;
			{8'd19, 8'd80}: color_data = 12'hba8;
			{8'd19, 8'd81}: color_data = 12'hfec;
			{8'd19, 8'd82}: color_data = 12'hfec;
			{8'd19, 8'd83}: color_data = 12'hfeb;
			{8'd19, 8'd84}: color_data = 12'hfeb;
			{8'd19, 8'd85}: color_data = 12'hfdb;
			{8'd19, 8'd86}: color_data = 12'h765;
			{8'd19, 8'd87}: color_data = 12'h000;
			{8'd19, 8'd97}: color_data = 12'h010;
			{8'd19, 8'd98}: color_data = 12'h072;
			{8'd19, 8'd99}: color_data = 12'h093;
			{8'd19, 8'd100}: color_data = 12'h374;
			{8'd19, 8'd101}: color_data = 12'h8a9;
			{8'd19, 8'd102}: color_data = 12'hddd;
			{8'd19, 8'd103}: color_data = 12'hfff;
			{8'd19, 8'd104}: color_data = 12'hfff;
			{8'd19, 8'd105}: color_data = 12'hfff;
			{8'd19, 8'd106}: color_data = 12'heee;
			{8'd19, 8'd107}: color_data = 12'h999;
			{8'd19, 8'd108}: color_data = 12'h111;
			{8'd19, 8'd109}: color_data = 12'h000;
			{8'd19, 8'd110}: color_data = 12'h011;
			{8'd19, 8'd111}: color_data = 12'h013;
			{8'd19, 8'd112}: color_data = 12'h013;
			{8'd19, 8'd113}: color_data = 12'h124;
			{8'd19, 8'd114}: color_data = 12'h124;
			{8'd19, 8'd115}: color_data = 12'h124;
			{8'd19, 8'd116}: color_data = 12'h124;
			{8'd19, 8'd117}: color_data = 12'h123;
			{8'd19, 8'd118}: color_data = 12'h012;
			{8'd19, 8'd119}: color_data = 12'h000;
			{8'd19, 8'd120}: color_data = 12'h000;
			{8'd19, 8'd127}: color_data = 12'h000;
			{8'd19, 8'd128}: color_data = 12'h001;
			{8'd19, 8'd129}: color_data = 12'h013;
			{8'd19, 8'd130}: color_data = 12'h125;
			{8'd19, 8'd131}: color_data = 12'h136;
			{8'd19, 8'd132}: color_data = 12'h247;
			{8'd19, 8'd133}: color_data = 12'h247;
			{8'd19, 8'd134}: color_data = 12'h136;
			{8'd19, 8'd135}: color_data = 12'h012;
			{8'd19, 8'd137}: color_data = 12'h000;
			{8'd19, 8'd138}: color_data = 12'h532;
			{8'd19, 8'd139}: color_data = 12'h643;
			{8'd19, 8'd140}: color_data = 12'h633;
			{8'd19, 8'd141}: color_data = 12'h633;
			{8'd19, 8'd142}: color_data = 12'h633;
			{8'd19, 8'd143}: color_data = 12'h633;
			{8'd19, 8'd144}: color_data = 12'h633;
			{8'd19, 8'd145}: color_data = 12'h653;
			{8'd19, 8'd146}: color_data = 12'h543;
			{8'd20, 8'd20}: color_data = 12'hfc5;
			{8'd20, 8'd21}: color_data = 12'hfc5;
			{8'd20, 8'd22}: color_data = 12'heb2;
			{8'd20, 8'd23}: color_data = 12'hd90;
			{8'd20, 8'd24}: color_data = 12'hd90;
			{8'd20, 8'd25}: color_data = 12'hd90;
			{8'd20, 8'd26}: color_data = 12'hd90;
			{8'd20, 8'd27}: color_data = 12'hd90;
			{8'd20, 8'd28}: color_data = 12'hd90;
			{8'd20, 8'd29}: color_data = 12'hd90;
			{8'd20, 8'd30}: color_data = 12'hd90;
			{8'd20, 8'd31}: color_data = 12'hd90;
			{8'd20, 8'd32}: color_data = 12'hd90;
			{8'd20, 8'd33}: color_data = 12'hd90;
			{8'd20, 8'd34}: color_data = 12'hd90;
			{8'd20, 8'd35}: color_data = 12'hd90;
			{8'd20, 8'd36}: color_data = 12'heb2;
			{8'd20, 8'd37}: color_data = 12'hfc5;
			{8'd20, 8'd38}: color_data = 12'hfc5;
			{8'd20, 8'd56}: color_data = 12'h000;
			{8'd20, 8'd57}: color_data = 12'h041;
			{8'd20, 8'd58}: color_data = 12'h083;
			{8'd20, 8'd59}: color_data = 12'h0a4;
			{8'd20, 8'd60}: color_data = 12'h0a3;
			{8'd20, 8'd61}: color_data = 12'h0a3;
			{8'd20, 8'd62}: color_data = 12'h0a3;
			{8'd20, 8'd63}: color_data = 12'h0a3;
			{8'd20, 8'd64}: color_data = 12'h0a3;
			{8'd20, 8'd65}: color_data = 12'h0a3;
			{8'd20, 8'd66}: color_data = 12'h0a3;
			{8'd20, 8'd67}: color_data = 12'h0a3;
			{8'd20, 8'd68}: color_data = 12'h0a3;
			{8'd20, 8'd69}: color_data = 12'h0a3;
			{8'd20, 8'd70}: color_data = 12'h0a3;
			{8'd20, 8'd71}: color_data = 12'h0a3;
			{8'd20, 8'd72}: color_data = 12'h0a3;
			{8'd20, 8'd73}: color_data = 12'h0a3;
			{8'd20, 8'd74}: color_data = 12'h0a3;
			{8'd20, 8'd75}: color_data = 12'h0a3;
			{8'd20, 8'd76}: color_data = 12'h0a3;
			{8'd20, 8'd77}: color_data = 12'h241;
			{8'd20, 8'd78}: color_data = 12'h742;
			{8'd20, 8'd79}: color_data = 12'h643;
			{8'd20, 8'd80}: color_data = 12'hfdb;
			{8'd20, 8'd81}: color_data = 12'hfdb;
			{8'd20, 8'd82}: color_data = 12'hba8;
			{8'd20, 8'd83}: color_data = 12'hfda;
			{8'd20, 8'd84}: color_data = 12'hfdb;
			{8'd20, 8'd85}: color_data = 12'hfdb;
			{8'd20, 8'd86}: color_data = 12'hfdb;
			{8'd20, 8'd87}: color_data = 12'h876;
			{8'd20, 8'd88}: color_data = 12'h000;
			{8'd20, 8'd96}: color_data = 12'h000;
			{8'd20, 8'd97}: color_data = 12'h062;
			{8'd20, 8'd98}: color_data = 12'h051;
			{8'd20, 8'd99}: color_data = 12'h9a9;
			{8'd20, 8'd100}: color_data = 12'hfff;
			{8'd20, 8'd101}: color_data = 12'hfff;
			{8'd20, 8'd102}: color_data = 12'hddd;
			{8'd20, 8'd103}: color_data = 12'hbbb;
			{8'd20, 8'd104}: color_data = 12'hbbb;
			{8'd20, 8'd105}: color_data = 12'heee;
			{8'd20, 8'd106}: color_data = 12'hfff;
			{8'd20, 8'd107}: color_data = 12'hfff;
			{8'd20, 8'd108}: color_data = 12'h777;
			{8'd20, 8'd109}: color_data = 12'h125;
			{8'd20, 8'd110}: color_data = 12'h248;
			{8'd20, 8'd111}: color_data = 12'h249;
			{8'd20, 8'd112}: color_data = 12'h249;
			{8'd20, 8'd113}: color_data = 12'h249;
			{8'd20, 8'd114}: color_data = 12'h249;
			{8'd20, 8'd115}: color_data = 12'h249;
			{8'd20, 8'd116}: color_data = 12'h249;
			{8'd20, 8'd117}: color_data = 12'h249;
			{8'd20, 8'd118}: color_data = 12'h248;
			{8'd20, 8'd119}: color_data = 12'h137;
			{8'd20, 8'd120}: color_data = 12'h124;
			{8'd20, 8'd121}: color_data = 12'h001;
			{8'd20, 8'd125}: color_data = 12'h000;
			{8'd20, 8'd126}: color_data = 12'h012;
			{8'd20, 8'd127}: color_data = 12'h125;
			{8'd20, 8'd128}: color_data = 12'h247;
			{8'd20, 8'd129}: color_data = 12'h249;
			{8'd20, 8'd130}: color_data = 12'h249;
			{8'd20, 8'd131}: color_data = 12'h249;
			{8'd20, 8'd132}: color_data = 12'h249;
			{8'd20, 8'd133}: color_data = 12'h249;
			{8'd20, 8'd134}: color_data = 12'h259;
			{8'd20, 8'd135}: color_data = 12'h248;
			{8'd20, 8'd136}: color_data = 12'h013;
			{8'd20, 8'd137}: color_data = 12'h100;
			{8'd20, 8'd138}: color_data = 12'h633;
			{8'd20, 8'd139}: color_data = 12'h643;
			{8'd20, 8'd140}: color_data = 12'h633;
			{8'd20, 8'd141}: color_data = 12'h633;
			{8'd20, 8'd142}: color_data = 12'h633;
			{8'd20, 8'd143}: color_data = 12'h633;
			{8'd20, 8'd144}: color_data = 12'h633;
			{8'd20, 8'd145}: color_data = 12'h643;
			{8'd20, 8'd146}: color_data = 12'h542;
			{8'd21, 8'd20}: color_data = 12'hfc4;
			{8'd21, 8'd21}: color_data = 12'hfc5;
			{8'd21, 8'd22}: color_data = 12'hea1;
			{8'd21, 8'd23}: color_data = 12'hd90;
			{8'd21, 8'd24}: color_data = 12'hd90;
			{8'd21, 8'd25}: color_data = 12'hd90;
			{8'd21, 8'd26}: color_data = 12'hd90;
			{8'd21, 8'd27}: color_data = 12'hd90;
			{8'd21, 8'd28}: color_data = 12'hd90;
			{8'd21, 8'd29}: color_data = 12'hd90;
			{8'd21, 8'd30}: color_data = 12'hd90;
			{8'd21, 8'd31}: color_data = 12'hd90;
			{8'd21, 8'd32}: color_data = 12'hd90;
			{8'd21, 8'd33}: color_data = 12'hd90;
			{8'd21, 8'd34}: color_data = 12'hd90;
			{8'd21, 8'd35}: color_data = 12'hd90;
			{8'd21, 8'd36}: color_data = 12'heb2;
			{8'd21, 8'd37}: color_data = 12'hfc5;
			{8'd21, 8'd38}: color_data = 12'hfc4;
			{8'd21, 8'd55}: color_data = 12'h010;
			{8'd21, 8'd56}: color_data = 12'h062;
			{8'd21, 8'd57}: color_data = 12'h0a3;
			{8'd21, 8'd58}: color_data = 12'h0a3;
			{8'd21, 8'd59}: color_data = 12'h0a3;
			{8'd21, 8'd60}: color_data = 12'h0a3;
			{8'd21, 8'd61}: color_data = 12'h0a3;
			{8'd21, 8'd62}: color_data = 12'h0a3;
			{8'd21, 8'd63}: color_data = 12'h0a3;
			{8'd21, 8'd64}: color_data = 12'h0a3;
			{8'd21, 8'd65}: color_data = 12'h0a3;
			{8'd21, 8'd66}: color_data = 12'h0a3;
			{8'd21, 8'd67}: color_data = 12'h0a3;
			{8'd21, 8'd68}: color_data = 12'h0a3;
			{8'd21, 8'd69}: color_data = 12'h0a3;
			{8'd21, 8'd70}: color_data = 12'h0a3;
			{8'd21, 8'd71}: color_data = 12'h0a3;
			{8'd21, 8'd72}: color_data = 12'h0a3;
			{8'd21, 8'd73}: color_data = 12'h0a3;
			{8'd21, 8'd74}: color_data = 12'h0a3;
			{8'd21, 8'd75}: color_data = 12'h0a3;
			{8'd21, 8'd76}: color_data = 12'h142;
			{8'd21, 8'd77}: color_data = 12'h742;
			{8'd21, 8'd78}: color_data = 12'h842;
			{8'd21, 8'd79}: color_data = 12'h632;
			{8'd21, 8'd80}: color_data = 12'hcb9;
			{8'd21, 8'd81}: color_data = 12'hca8;
			{8'd21, 8'd82}: color_data = 12'hb98;
			{8'd21, 8'd83}: color_data = 12'heda;
			{8'd21, 8'd84}: color_data = 12'hca8;
			{8'd21, 8'd85}: color_data = 12'heca;
			{8'd21, 8'd86}: color_data = 12'hfdb;
			{8'd21, 8'd87}: color_data = 12'hfdb;
			{8'd21, 8'd88}: color_data = 12'h543;
			{8'd21, 8'd95}: color_data = 12'h000;
			{8'd21, 8'd96}: color_data = 12'h021;
			{8'd21, 8'd97}: color_data = 12'h183;
			{8'd21, 8'd98}: color_data = 12'h354;
			{8'd21, 8'd99}: color_data = 12'ha9a;
			{8'd21, 8'd100}: color_data = 12'h999;
			{8'd21, 8'd101}: color_data = 12'h888;
			{8'd21, 8'd102}: color_data = 12'h888;
			{8'd21, 8'd103}: color_data = 12'hbbb;
			{8'd21, 8'd104}: color_data = 12'hddd;
			{8'd21, 8'd105}: color_data = 12'hccc;
			{8'd21, 8'd106}: color_data = 12'hfff;
			{8'd21, 8'd107}: color_data = 12'heef;
			{8'd21, 8'd108}: color_data = 12'h457;
			{8'd21, 8'd109}: color_data = 12'h136;
			{8'd21, 8'd110}: color_data = 12'h135;
			{8'd21, 8'd111}: color_data = 12'h248;
			{8'd21, 8'd112}: color_data = 12'h249;
			{8'd21, 8'd113}: color_data = 12'h249;
			{8'd21, 8'd114}: color_data = 12'h249;
			{8'd21, 8'd115}: color_data = 12'h249;
			{8'd21, 8'd116}: color_data = 12'h249;
			{8'd21, 8'd117}: color_data = 12'h249;
			{8'd21, 8'd118}: color_data = 12'h249;
			{8'd21, 8'd119}: color_data = 12'h249;
			{8'd21, 8'd120}: color_data = 12'h249;
			{8'd21, 8'd121}: color_data = 12'h137;
			{8'd21, 8'd122}: color_data = 12'h013;
			{8'd21, 8'd123}: color_data = 12'h000;
			{8'd21, 8'd124}: color_data = 12'h001;
			{8'd21, 8'd125}: color_data = 12'h125;
			{8'd21, 8'd126}: color_data = 12'h248;
			{8'd21, 8'd127}: color_data = 12'h249;
			{8'd21, 8'd128}: color_data = 12'h249;
			{8'd21, 8'd129}: color_data = 12'h249;
			{8'd21, 8'd130}: color_data = 12'h249;
			{8'd21, 8'd131}: color_data = 12'h249;
			{8'd21, 8'd132}: color_data = 12'h249;
			{8'd21, 8'd133}: color_data = 12'h249;
			{8'd21, 8'd134}: color_data = 12'h249;
			{8'd21, 8'd135}: color_data = 12'h249;
			{8'd21, 8'd136}: color_data = 12'h147;
			{8'd21, 8'd137}: color_data = 12'h111;
			{8'd21, 8'd138}: color_data = 12'h633;
			{8'd21, 8'd139}: color_data = 12'h633;
			{8'd21, 8'd140}: color_data = 12'h633;
			{8'd21, 8'd141}: color_data = 12'h633;
			{8'd21, 8'd142}: color_data = 12'h633;
			{8'd21, 8'd143}: color_data = 12'h633;
			{8'd21, 8'd144}: color_data = 12'h633;
			{8'd21, 8'd145}: color_data = 12'h543;
			{8'd21, 8'd146}: color_data = 12'h432;
			{8'd22, 8'd19}: color_data = 12'hfb6;
			{8'd22, 8'd20}: color_data = 12'hfc5;
			{8'd22, 8'd21}: color_data = 12'hfc5;
			{8'd22, 8'd22}: color_data = 12'hea1;
			{8'd22, 8'd23}: color_data = 12'hd90;
			{8'd22, 8'd24}: color_data = 12'hd90;
			{8'd22, 8'd25}: color_data = 12'hd90;
			{8'd22, 8'd26}: color_data = 12'hea2;
			{8'd22, 8'd27}: color_data = 12'hfb3;
			{8'd22, 8'd28}: color_data = 12'hd90;
			{8'd22, 8'd29}: color_data = 12'hd90;
			{8'd22, 8'd30}: color_data = 12'hd90;
			{8'd22, 8'd31}: color_data = 12'hd90;
			{8'd22, 8'd32}: color_data = 12'hd90;
			{8'd22, 8'd33}: color_data = 12'hd90;
			{8'd22, 8'd34}: color_data = 12'hd90;
			{8'd22, 8'd35}: color_data = 12'hd90;
			{8'd22, 8'd36}: color_data = 12'hfc4;
			{8'd22, 8'd37}: color_data = 12'hfc5;
			{8'd22, 8'd38}: color_data = 12'hfc5;
			{8'd22, 8'd54}: color_data = 12'h020;
			{8'd22, 8'd55}: color_data = 12'h082;
			{8'd22, 8'd56}: color_data = 12'h0a4;
			{8'd22, 8'd57}: color_data = 12'h0a3;
			{8'd22, 8'd58}: color_data = 12'h0a3;
			{8'd22, 8'd59}: color_data = 12'h0a3;
			{8'd22, 8'd60}: color_data = 12'h0a3;
			{8'd22, 8'd61}: color_data = 12'h0a3;
			{8'd22, 8'd62}: color_data = 12'h0a3;
			{8'd22, 8'd63}: color_data = 12'h0a3;
			{8'd22, 8'd64}: color_data = 12'h0a3;
			{8'd22, 8'd65}: color_data = 12'h0a3;
			{8'd22, 8'd66}: color_data = 12'h0a3;
			{8'd22, 8'd67}: color_data = 12'h0a3;
			{8'd22, 8'd68}: color_data = 12'h0a3;
			{8'd22, 8'd69}: color_data = 12'h0a3;
			{8'd22, 8'd70}: color_data = 12'h0a3;
			{8'd22, 8'd71}: color_data = 12'h0a3;
			{8'd22, 8'd72}: color_data = 12'h0a3;
			{8'd22, 8'd73}: color_data = 12'h0a3;
			{8'd22, 8'd74}: color_data = 12'h0a3;
			{8'd22, 8'd75}: color_data = 12'h152;
			{8'd22, 8'd76}: color_data = 12'h732;
			{8'd22, 8'd77}: color_data = 12'h842;
			{8'd22, 8'd78}: color_data = 12'h842;
			{8'd22, 8'd79}: color_data = 12'h842;
			{8'd22, 8'd80}: color_data = 12'h643;
			{8'd22, 8'd81}: color_data = 12'hdb9;
			{8'd22, 8'd82}: color_data = 12'ha87;
			{8'd22, 8'd83}: color_data = 12'h986;
			{8'd22, 8'd84}: color_data = 12'hca8;
			{8'd22, 8'd85}: color_data = 12'hdb9;
			{8'd22, 8'd86}: color_data = 12'hfdb;
			{8'd22, 8'd87}: color_data = 12'hfeb;
			{8'd22, 8'd88}: color_data = 12'h876;
			{8'd22, 8'd89}: color_data = 12'h000;
			{8'd22, 8'd90}: color_data = 12'h000;
			{8'd22, 8'd95}: color_data = 12'h222;
			{8'd22, 8'd96}: color_data = 12'haaa;
			{8'd22, 8'd97}: color_data = 12'hfef;
			{8'd22, 8'd98}: color_data = 12'hfff;
			{8'd22, 8'd99}: color_data = 12'hfff;
			{8'd22, 8'd100}: color_data = 12'hccc;
			{8'd22, 8'd101}: color_data = 12'heee;
			{8'd22, 8'd102}: color_data = 12'hccc;
			{8'd22, 8'd103}: color_data = 12'hccc;
			{8'd22, 8'd104}: color_data = 12'hfff;
			{8'd22, 8'd105}: color_data = 12'hfff;
			{8'd22, 8'd106}: color_data = 12'hbbb;
			{8'd22, 8'd107}: color_data = 12'h773;
			{8'd22, 8'd108}: color_data = 12'h136;
			{8'd22, 8'd109}: color_data = 12'h259;
			{8'd22, 8'd110}: color_data = 12'h237;
			{8'd22, 8'd111}: color_data = 12'h136;
			{8'd22, 8'd112}: color_data = 12'h249;
			{8'd22, 8'd113}: color_data = 12'h249;
			{8'd22, 8'd114}: color_data = 12'h249;
			{8'd22, 8'd115}: color_data = 12'h249;
			{8'd22, 8'd116}: color_data = 12'h249;
			{8'd22, 8'd117}: color_data = 12'h249;
			{8'd22, 8'd118}: color_data = 12'h249;
			{8'd22, 8'd119}: color_data = 12'h249;
			{8'd22, 8'd120}: color_data = 12'h249;
			{8'd22, 8'd121}: color_data = 12'h249;
			{8'd22, 8'd122}: color_data = 12'h248;
			{8'd22, 8'd123}: color_data = 12'h125;
			{8'd22, 8'd124}: color_data = 12'h247;
			{8'd22, 8'd125}: color_data = 12'h249;
			{8'd22, 8'd126}: color_data = 12'h249;
			{8'd22, 8'd127}: color_data = 12'h249;
			{8'd22, 8'd128}: color_data = 12'h249;
			{8'd22, 8'd129}: color_data = 12'h249;
			{8'd22, 8'd130}: color_data = 12'h249;
			{8'd22, 8'd131}: color_data = 12'h249;
			{8'd22, 8'd132}: color_data = 12'h249;
			{8'd22, 8'd133}: color_data = 12'h249;
			{8'd22, 8'd134}: color_data = 12'h249;
			{8'd22, 8'd135}: color_data = 12'h249;
			{8'd22, 8'd136}: color_data = 12'h249;
			{8'd22, 8'd137}: color_data = 12'h224;
			{8'd22, 8'd138}: color_data = 12'h633;
			{8'd22, 8'd139}: color_data = 12'h633;
			{8'd22, 8'd140}: color_data = 12'h633;
			{8'd22, 8'd141}: color_data = 12'h633;
			{8'd22, 8'd142}: color_data = 12'h633;
			{8'd22, 8'd143}: color_data = 12'h633;
			{8'd22, 8'd144}: color_data = 12'h633;
			{8'd22, 8'd145}: color_data = 12'h532;
			{8'd22, 8'd146}: color_data = 12'h331;
			{8'd23, 8'd19}: color_data = 12'hfc5;
			{8'd23, 8'd20}: color_data = 12'hfc5;
			{8'd23, 8'd21}: color_data = 12'hfc4;
			{8'd23, 8'd22}: color_data = 12'hda0;
			{8'd23, 8'd23}: color_data = 12'hd90;
			{8'd23, 8'd24}: color_data = 12'hd90;
			{8'd23, 8'd25}: color_data = 12'hd90;
			{8'd23, 8'd26}: color_data = 12'hfc4;
			{8'd23, 8'd27}: color_data = 12'hfb3;
			{8'd23, 8'd28}: color_data = 12'hd90;
			{8'd23, 8'd29}: color_data = 12'hd90;
			{8'd23, 8'd30}: color_data = 12'hd90;
			{8'd23, 8'd31}: color_data = 12'heb2;
			{8'd23, 8'd32}: color_data = 12'hd90;
			{8'd23, 8'd33}: color_data = 12'hd90;
			{8'd23, 8'd34}: color_data = 12'hd90;
			{8'd23, 8'd35}: color_data = 12'hda0;
			{8'd23, 8'd36}: color_data = 12'hfc4;
			{8'd23, 8'd37}: color_data = 12'hfc4;
			{8'd23, 8'd38}: color_data = 12'hfc5;
			{8'd23, 8'd53}: color_data = 12'h020;
			{8'd23, 8'd54}: color_data = 12'h083;
			{8'd23, 8'd55}: color_data = 12'h0a3;
			{8'd23, 8'd56}: color_data = 12'h0a3;
			{8'd23, 8'd57}: color_data = 12'h0a3;
			{8'd23, 8'd58}: color_data = 12'h0a3;
			{8'd23, 8'd59}: color_data = 12'h0a3;
			{8'd23, 8'd60}: color_data = 12'h0a3;
			{8'd23, 8'd61}: color_data = 12'h0a3;
			{8'd23, 8'd62}: color_data = 12'h0a3;
			{8'd23, 8'd63}: color_data = 12'h0a3;
			{8'd23, 8'd64}: color_data = 12'h0a3;
			{8'd23, 8'd65}: color_data = 12'h0a3;
			{8'd23, 8'd66}: color_data = 12'h0a3;
			{8'd23, 8'd67}: color_data = 12'h0a3;
			{8'd23, 8'd68}: color_data = 12'h0a3;
			{8'd23, 8'd69}: color_data = 12'h0a3;
			{8'd23, 8'd70}: color_data = 12'h0a3;
			{8'd23, 8'd71}: color_data = 12'h0a3;
			{8'd23, 8'd72}: color_data = 12'h0a3;
			{8'd23, 8'd73}: color_data = 12'h0a3;
			{8'd23, 8'd74}: color_data = 12'h152;
			{8'd23, 8'd75}: color_data = 12'h732;
			{8'd23, 8'd76}: color_data = 12'h842;
			{8'd23, 8'd77}: color_data = 12'h631;
			{8'd23, 8'd78}: color_data = 12'h842;
			{8'd23, 8'd79}: color_data = 12'h842;
			{8'd23, 8'd80}: color_data = 12'h742;
			{8'd23, 8'd81}: color_data = 12'h643;
			{8'd23, 8'd82}: color_data = 12'hba8;
			{8'd23, 8'd83}: color_data = 12'h876;
			{8'd23, 8'd84}: color_data = 12'heca;
			{8'd23, 8'd85}: color_data = 12'hfeb;
			{8'd23, 8'd86}: color_data = 12'hfdb;
			{8'd23, 8'd87}: color_data = 12'hfeb;
			{8'd23, 8'd88}: color_data = 12'h665;
			{8'd23, 8'd89}: color_data = 12'h310;
			{8'd23, 8'd90}: color_data = 12'h321;
			{8'd23, 8'd94}: color_data = 12'h000;
			{8'd23, 8'd95}: color_data = 12'h455;
			{8'd23, 8'd96}: color_data = 12'hfff;
			{8'd23, 8'd97}: color_data = 12'hfff;
			{8'd23, 8'd98}: color_data = 12'hfff;
			{8'd23, 8'd99}: color_data = 12'hfff;
			{8'd23, 8'd100}: color_data = 12'hfff;
			{8'd23, 8'd101}: color_data = 12'hfff;
			{8'd23, 8'd102}: color_data = 12'hfff;
			{8'd23, 8'd103}: color_data = 12'hfff;
			{8'd23, 8'd104}: color_data = 12'hfff;
			{8'd23, 8'd105}: color_data = 12'heee;
			{8'd23, 8'd106}: color_data = 12'h881;
			{8'd23, 8'd107}: color_data = 12'hff0;
			{8'd23, 8'd108}: color_data = 12'h553;
			{8'd23, 8'd109}: color_data = 12'h249;
			{8'd23, 8'd110}: color_data = 12'h248;
			{8'd23, 8'd111}: color_data = 12'h135;
			{8'd23, 8'd112}: color_data = 12'h249;
			{8'd23, 8'd113}: color_data = 12'h249;
			{8'd23, 8'd114}: color_data = 12'h249;
			{8'd23, 8'd115}: color_data = 12'h249;
			{8'd23, 8'd116}: color_data = 12'h249;
			{8'd23, 8'd117}: color_data = 12'h249;
			{8'd23, 8'd118}: color_data = 12'h249;
			{8'd23, 8'd119}: color_data = 12'h249;
			{8'd23, 8'd120}: color_data = 12'h249;
			{8'd23, 8'd121}: color_data = 12'h249;
			{8'd23, 8'd122}: color_data = 12'h249;
			{8'd23, 8'd123}: color_data = 12'h249;
			{8'd23, 8'd124}: color_data = 12'h249;
			{8'd23, 8'd125}: color_data = 12'h249;
			{8'd23, 8'd126}: color_data = 12'h249;
			{8'd23, 8'd127}: color_data = 12'h249;
			{8'd23, 8'd128}: color_data = 12'h249;
			{8'd23, 8'd129}: color_data = 12'h249;
			{8'd23, 8'd130}: color_data = 12'h249;
			{8'd23, 8'd131}: color_data = 12'h249;
			{8'd23, 8'd132}: color_data = 12'h249;
			{8'd23, 8'd133}: color_data = 12'h249;
			{8'd23, 8'd134}: color_data = 12'h249;
			{8'd23, 8'd135}: color_data = 12'h249;
			{8'd23, 8'd136}: color_data = 12'h249;
			{8'd23, 8'd137}: color_data = 12'h125;
			{8'd23, 8'd138}: color_data = 12'h422;
			{8'd23, 8'd139}: color_data = 12'h643;
			{8'd23, 8'd140}: color_data = 12'h633;
			{8'd23, 8'd141}: color_data = 12'h633;
			{8'd23, 8'd142}: color_data = 12'h633;
			{8'd23, 8'd143}: color_data = 12'h633;
			{8'd23, 8'd144}: color_data = 12'h633;
			{8'd23, 8'd145}: color_data = 12'h542;
			{8'd23, 8'd146}: color_data = 12'h221;
			{8'd24, 8'd19}: color_data = 12'hfc5;
			{8'd24, 8'd20}: color_data = 12'hfc4;
			{8'd24, 8'd21}: color_data = 12'hfb3;
			{8'd24, 8'd22}: color_data = 12'hd90;
			{8'd24, 8'd23}: color_data = 12'hd90;
			{8'd24, 8'd24}: color_data = 12'hd90;
			{8'd24, 8'd25}: color_data = 12'hda0;
			{8'd24, 8'd26}: color_data = 12'hfc6;
			{8'd24, 8'd27}: color_data = 12'heb2;
			{8'd24, 8'd28}: color_data = 12'hd90;
			{8'd24, 8'd29}: color_data = 12'hd90;
			{8'd24, 8'd30}: color_data = 12'hea1;
			{8'd24, 8'd31}: color_data = 12'hfc5;
			{8'd24, 8'd32}: color_data = 12'hea0;
			{8'd24, 8'd33}: color_data = 12'hd90;
			{8'd24, 8'd34}: color_data = 12'hd90;
			{8'd24, 8'd35}: color_data = 12'hea1;
			{8'd24, 8'd36}: color_data = 12'hfc5;
			{8'd24, 8'd37}: color_data = 12'hfc5;
			{8'd24, 8'd38}: color_data = 12'hff7;
			{8'd24, 8'd52}: color_data = 12'h010;
			{8'd24, 8'd53}: color_data = 12'h082;
			{8'd24, 8'd54}: color_data = 12'h0a3;
			{8'd24, 8'd55}: color_data = 12'h0a3;
			{8'd24, 8'd56}: color_data = 12'h0a3;
			{8'd24, 8'd57}: color_data = 12'h0a3;
			{8'd24, 8'd58}: color_data = 12'h0a3;
			{8'd24, 8'd59}: color_data = 12'h0a3;
			{8'd24, 8'd60}: color_data = 12'h0a3;
			{8'd24, 8'd61}: color_data = 12'h0a3;
			{8'd24, 8'd62}: color_data = 12'h0a3;
			{8'd24, 8'd63}: color_data = 12'h0a3;
			{8'd24, 8'd64}: color_data = 12'h0a3;
			{8'd24, 8'd65}: color_data = 12'h0a3;
			{8'd24, 8'd66}: color_data = 12'h0a3;
			{8'd24, 8'd67}: color_data = 12'h0a3;
			{8'd24, 8'd68}: color_data = 12'h0a3;
			{8'd24, 8'd69}: color_data = 12'h0a3;
			{8'd24, 8'd70}: color_data = 12'h0a3;
			{8'd24, 8'd71}: color_data = 12'h0a3;
			{8'd24, 8'd72}: color_data = 12'h0a3;
			{8'd24, 8'd73}: color_data = 12'h051;
			{8'd24, 8'd74}: color_data = 12'h631;
			{8'd24, 8'd75}: color_data = 12'h741;
			{8'd24, 8'd76}: color_data = 12'h632;
			{8'd24, 8'd77}: color_data = 12'h986;
			{8'd24, 8'd78}: color_data = 12'h642;
			{8'd24, 8'd79}: color_data = 12'h842;
			{8'd24, 8'd80}: color_data = 12'h842;
			{8'd24, 8'd81}: color_data = 12'h742;
			{8'd24, 8'd82}: color_data = 12'h643;
			{8'd24, 8'd83}: color_data = 12'hb98;
			{8'd24, 8'd84}: color_data = 12'h987;
			{8'd24, 8'd85}: color_data = 12'hdb9;
			{8'd24, 8'd86}: color_data = 12'hfdb;
			{8'd24, 8'd87}: color_data = 12'heda;
			{8'd24, 8'd88}: color_data = 12'h542;
			{8'd24, 8'd89}: color_data = 12'h842;
			{8'd24, 8'd90}: color_data = 12'h321;
			{8'd24, 8'd93}: color_data = 12'h000;
			{8'd24, 8'd94}: color_data = 12'h041;
			{8'd24, 8'd95}: color_data = 12'h485;
			{8'd24, 8'd96}: color_data = 12'hfff;
			{8'd24, 8'd97}: color_data = 12'hfff;
			{8'd24, 8'd98}: color_data = 12'hfff;
			{8'd24, 8'd99}: color_data = 12'hfff;
			{8'd24, 8'd100}: color_data = 12'hfff;
			{8'd24, 8'd101}: color_data = 12'hfff;
			{8'd24, 8'd102}: color_data = 12'hfff;
			{8'd24, 8'd103}: color_data = 12'hfff;
			{8'd24, 8'd104}: color_data = 12'hfff;
			{8'd24, 8'd105}: color_data = 12'hfff;
			{8'd24, 8'd106}: color_data = 12'h983;
			{8'd24, 8'd107}: color_data = 12'h990;
			{8'd24, 8'd108}: color_data = 12'h236;
			{8'd24, 8'd109}: color_data = 12'h137;
			{8'd24, 8'd110}: color_data = 12'h125;
			{8'd24, 8'd111}: color_data = 12'h248;
			{8'd24, 8'd112}: color_data = 12'h249;
			{8'd24, 8'd113}: color_data = 12'h249;
			{8'd24, 8'd114}: color_data = 12'h249;
			{8'd24, 8'd115}: color_data = 12'h249;
			{8'd24, 8'd116}: color_data = 12'h249;
			{8'd24, 8'd117}: color_data = 12'h249;
			{8'd24, 8'd118}: color_data = 12'h249;
			{8'd24, 8'd119}: color_data = 12'h249;
			{8'd24, 8'd120}: color_data = 12'h249;
			{8'd24, 8'd121}: color_data = 12'h249;
			{8'd24, 8'd122}: color_data = 12'h249;
			{8'd24, 8'd123}: color_data = 12'h249;
			{8'd24, 8'd124}: color_data = 12'h249;
			{8'd24, 8'd125}: color_data = 12'h249;
			{8'd24, 8'd126}: color_data = 12'h249;
			{8'd24, 8'd127}: color_data = 12'h249;
			{8'd24, 8'd128}: color_data = 12'h249;
			{8'd24, 8'd129}: color_data = 12'h249;
			{8'd24, 8'd130}: color_data = 12'h249;
			{8'd24, 8'd131}: color_data = 12'h249;
			{8'd24, 8'd132}: color_data = 12'h249;
			{8'd24, 8'd133}: color_data = 12'h249;
			{8'd24, 8'd134}: color_data = 12'h249;
			{8'd24, 8'd135}: color_data = 12'h249;
			{8'd24, 8'd136}: color_data = 12'h249;
			{8'd24, 8'd137}: color_data = 12'h137;
			{8'd24, 8'd138}: color_data = 12'h112;
			{8'd24, 8'd139}: color_data = 12'h422;
			{8'd24, 8'd140}: color_data = 12'h633;
			{8'd24, 8'd141}: color_data = 12'h633;
			{8'd24, 8'd142}: color_data = 12'h633;
			{8'd24, 8'd143}: color_data = 12'h643;
			{8'd24, 8'd144}: color_data = 12'h532;
			{8'd24, 8'd145}: color_data = 12'h542;
			{8'd24, 8'd146}: color_data = 12'h000;
			{8'd25, 8'd19}: color_data = 12'hfc5;
			{8'd25, 8'd20}: color_data = 12'hfc5;
			{8'd25, 8'd21}: color_data = 12'heb2;
			{8'd25, 8'd22}: color_data = 12'hd90;
			{8'd25, 8'd23}: color_data = 12'hd90;
			{8'd25, 8'd24}: color_data = 12'hd90;
			{8'd25, 8'd25}: color_data = 12'heb2;
			{8'd25, 8'd26}: color_data = 12'hfd7;
			{8'd25, 8'd27}: color_data = 12'hea1;
			{8'd25, 8'd28}: color_data = 12'hd90;
			{8'd25, 8'd29}: color_data = 12'hd90;
			{8'd25, 8'd30}: color_data = 12'heb2;
			{8'd25, 8'd31}: color_data = 12'hfc5;
			{8'd25, 8'd32}: color_data = 12'hd90;
			{8'd25, 8'd33}: color_data = 12'hd90;
			{8'd25, 8'd34}: color_data = 12'hd90;
			{8'd25, 8'd35}: color_data = 12'heb2;
			{8'd25, 8'd36}: color_data = 12'hfc5;
			{8'd25, 8'd37}: color_data = 12'hfc5;
			{8'd25, 8'd51}: color_data = 12'h000;
			{8'd25, 8'd52}: color_data = 12'h062;
			{8'd25, 8'd53}: color_data = 12'h0a4;
			{8'd25, 8'd54}: color_data = 12'h0a3;
			{8'd25, 8'd55}: color_data = 12'h0a3;
			{8'd25, 8'd56}: color_data = 12'h0a3;
			{8'd25, 8'd57}: color_data = 12'h0a3;
			{8'd25, 8'd58}: color_data = 12'h0a3;
			{8'd25, 8'd59}: color_data = 12'h0a3;
			{8'd25, 8'd60}: color_data = 12'h0a3;
			{8'd25, 8'd61}: color_data = 12'h0a3;
			{8'd25, 8'd62}: color_data = 12'h0a3;
			{8'd25, 8'd63}: color_data = 12'h0a3;
			{8'd25, 8'd64}: color_data = 12'h0a3;
			{8'd25, 8'd65}: color_data = 12'h0a3;
			{8'd25, 8'd66}: color_data = 12'h0a3;
			{8'd25, 8'd67}: color_data = 12'h0a3;
			{8'd25, 8'd68}: color_data = 12'h0a3;
			{8'd25, 8'd69}: color_data = 12'h0a3;
			{8'd25, 8'd70}: color_data = 12'h0a3;
			{8'd25, 8'd71}: color_data = 12'h093;
			{8'd25, 8'd72}: color_data = 12'h062;
			{8'd25, 8'd73}: color_data = 12'h121;
			{8'd25, 8'd74}: color_data = 12'h865;
			{8'd25, 8'd75}: color_data = 12'h986;
			{8'd25, 8'd76}: color_data = 12'hdb9;
			{8'd25, 8'd77}: color_data = 12'hfeb;
			{8'd25, 8'd78}: color_data = 12'h754;
			{8'd25, 8'd79}: color_data = 12'h842;
			{8'd25, 8'd80}: color_data = 12'h842;
			{8'd25, 8'd81}: color_data = 12'h842;
			{8'd25, 8'd82}: color_data = 12'h731;
			{8'd25, 8'd83}: color_data = 12'h865;
			{8'd25, 8'd84}: color_data = 12'hfdb;
			{8'd25, 8'd85}: color_data = 12'heca;
			{8'd25, 8'd86}: color_data = 12'hfdb;
			{8'd25, 8'd87}: color_data = 12'h976;
			{8'd25, 8'd88}: color_data = 12'h732;
			{8'd25, 8'd89}: color_data = 12'h842;
			{8'd25, 8'd90}: color_data = 12'h421;
			{8'd25, 8'd91}: color_data = 12'h000;
			{8'd25, 8'd93}: color_data = 12'h010;
			{8'd25, 8'd94}: color_data = 12'h062;
			{8'd25, 8'd95}: color_data = 12'h244;
			{8'd25, 8'd96}: color_data = 12'heee;
			{8'd25, 8'd97}: color_data = 12'hfff;
			{8'd25, 8'd98}: color_data = 12'hfff;
			{8'd25, 8'd99}: color_data = 12'hfff;
			{8'd25, 8'd100}: color_data = 12'hfff;
			{8'd25, 8'd101}: color_data = 12'hfff;
			{8'd25, 8'd102}: color_data = 12'hfff;
			{8'd25, 8'd103}: color_data = 12'hfff;
			{8'd25, 8'd104}: color_data = 12'hfff;
			{8'd25, 8'd105}: color_data = 12'hddd;
			{8'd25, 8'd106}: color_data = 12'h124;
			{8'd25, 8'd107}: color_data = 12'h025;
			{8'd25, 8'd108}: color_data = 12'h136;
			{8'd25, 8'd109}: color_data = 12'h137;
			{8'd25, 8'd110}: color_data = 12'h249;
			{8'd25, 8'd111}: color_data = 12'h249;
			{8'd25, 8'd112}: color_data = 12'h249;
			{8'd25, 8'd113}: color_data = 12'h249;
			{8'd25, 8'd114}: color_data = 12'h249;
			{8'd25, 8'd115}: color_data = 12'h249;
			{8'd25, 8'd116}: color_data = 12'h249;
			{8'd25, 8'd117}: color_data = 12'h249;
			{8'd25, 8'd118}: color_data = 12'h249;
			{8'd25, 8'd119}: color_data = 12'h249;
			{8'd25, 8'd120}: color_data = 12'h249;
			{8'd25, 8'd121}: color_data = 12'h249;
			{8'd25, 8'd122}: color_data = 12'h249;
			{8'd25, 8'd123}: color_data = 12'h249;
			{8'd25, 8'd124}: color_data = 12'h249;
			{8'd25, 8'd125}: color_data = 12'h249;
			{8'd25, 8'd126}: color_data = 12'h249;
			{8'd25, 8'd127}: color_data = 12'h249;
			{8'd25, 8'd128}: color_data = 12'h249;
			{8'd25, 8'd129}: color_data = 12'h249;
			{8'd25, 8'd130}: color_data = 12'h249;
			{8'd25, 8'd131}: color_data = 12'h249;
			{8'd25, 8'd132}: color_data = 12'h249;
			{8'd25, 8'd133}: color_data = 12'h249;
			{8'd25, 8'd134}: color_data = 12'h249;
			{8'd25, 8'd135}: color_data = 12'h249;
			{8'd25, 8'd136}: color_data = 12'h249;
			{8'd25, 8'd137}: color_data = 12'h249;
			{8'd25, 8'd138}: color_data = 12'h224;
			{8'd25, 8'd139}: color_data = 12'h532;
			{8'd25, 8'd140}: color_data = 12'h633;
			{8'd25, 8'd141}: color_data = 12'h633;
			{8'd25, 8'd142}: color_data = 12'h633;
			{8'd25, 8'd143}: color_data = 12'h633;
			{8'd25, 8'd144}: color_data = 12'h542;
			{8'd25, 8'd145}: color_data = 12'h542;
			{8'd26, 8'd19}: color_data = 12'hfc5;
			{8'd26, 8'd20}: color_data = 12'hfc5;
			{8'd26, 8'd21}: color_data = 12'hfc4;
			{8'd26, 8'd22}: color_data = 12'hfb3;
			{8'd26, 8'd23}: color_data = 12'hfb4;
			{8'd26, 8'd24}: color_data = 12'hfb3;
			{8'd26, 8'd25}: color_data = 12'hfc6;
			{8'd26, 8'd26}: color_data = 12'hfc5;
			{8'd26, 8'd27}: color_data = 12'hfc4;
			{8'd26, 8'd28}: color_data = 12'heb3;
			{8'd26, 8'd29}: color_data = 12'heb2;
			{8'd26, 8'd30}: color_data = 12'hfc5;
			{8'd26, 8'd31}: color_data = 12'hfb3;
			{8'd26, 8'd32}: color_data = 12'hd90;
			{8'd26, 8'd33}: color_data = 12'hd90;
			{8'd26, 8'd34}: color_data = 12'hd90;
			{8'd26, 8'd35}: color_data = 12'hfb3;
			{8'd26, 8'd36}: color_data = 12'hfc5;
			{8'd26, 8'd37}: color_data = 12'hfc5;
			{8'd26, 8'd51}: color_data = 12'h031;
			{8'd26, 8'd52}: color_data = 12'h0a3;
			{8'd26, 8'd53}: color_data = 12'h0a3;
			{8'd26, 8'd54}: color_data = 12'h0a3;
			{8'd26, 8'd55}: color_data = 12'h0a3;
			{8'd26, 8'd56}: color_data = 12'h0a3;
			{8'd26, 8'd57}: color_data = 12'h0a3;
			{8'd26, 8'd58}: color_data = 12'h0a3;
			{8'd26, 8'd59}: color_data = 12'h0a3;
			{8'd26, 8'd60}: color_data = 12'h0a3;
			{8'd26, 8'd61}: color_data = 12'h0a3;
			{8'd26, 8'd62}: color_data = 12'h0a3;
			{8'd26, 8'd63}: color_data = 12'h0a3;
			{8'd26, 8'd64}: color_data = 12'h0a3;
			{8'd26, 8'd65}: color_data = 12'h0a3;
			{8'd26, 8'd66}: color_data = 12'h0a3;
			{8'd26, 8'd67}: color_data = 12'h0a3;
			{8'd26, 8'd68}: color_data = 12'h0a3;
			{8'd26, 8'd69}: color_data = 12'h0a3;
			{8'd26, 8'd70}: color_data = 12'h093;
			{8'd26, 8'd71}: color_data = 12'h062;
			{8'd26, 8'd72}: color_data = 12'h093;
			{8'd26, 8'd73}: color_data = 12'h453;
			{8'd26, 8'd74}: color_data = 12'hfdb;
			{8'd26, 8'd75}: color_data = 12'hfeb;
			{8'd26, 8'd76}: color_data = 12'hfdb;
			{8'd26, 8'd77}: color_data = 12'hfdb;
			{8'd26, 8'd78}: color_data = 12'h865;
			{8'd26, 8'd79}: color_data = 12'h742;
			{8'd26, 8'd80}: color_data = 12'h631;
			{8'd26, 8'd81}: color_data = 12'h742;
			{8'd26, 8'd82}: color_data = 12'h531;
			{8'd26, 8'd83}: color_data = 12'hca9;
			{8'd26, 8'd84}: color_data = 12'hfdb;
			{8'd26, 8'd85}: color_data = 12'hfdb;
			{8'd26, 8'd86}: color_data = 12'hdca;
			{8'd26, 8'd87}: color_data = 12'h532;
			{8'd26, 8'd88}: color_data = 12'h842;
			{8'd26, 8'd89}: color_data = 12'h852;
			{8'd26, 8'd90}: color_data = 12'h421;
			{8'd26, 8'd91}: color_data = 12'h000;
			{8'd26, 8'd92}: color_data = 12'h000;
			{8'd26, 8'd93}: color_data = 12'h012;
			{8'd26, 8'd94}: color_data = 12'h247;
			{8'd26, 8'd95}: color_data = 12'h137;
			{8'd26, 8'd96}: color_data = 12'haab;
			{8'd26, 8'd97}: color_data = 12'hfff;
			{8'd26, 8'd98}: color_data = 12'hddd;
			{8'd26, 8'd99}: color_data = 12'heee;
			{8'd26, 8'd100}: color_data = 12'hfff;
			{8'd26, 8'd101}: color_data = 12'hfff;
			{8'd26, 8'd102}: color_data = 12'hccc;
			{8'd26, 8'd103}: color_data = 12'hbbb;
			{8'd26, 8'd104}: color_data = 12'hccc;
			{8'd26, 8'd105}: color_data = 12'h346;
			{8'd26, 8'd106}: color_data = 12'h136;
			{8'd26, 8'd107}: color_data = 12'h248;
			{8'd26, 8'd108}: color_data = 12'h249;
			{8'd26, 8'd109}: color_data = 12'h249;
			{8'd26, 8'd110}: color_data = 12'h249;
			{8'd26, 8'd111}: color_data = 12'h249;
			{8'd26, 8'd112}: color_data = 12'h249;
			{8'd26, 8'd113}: color_data = 12'h249;
			{8'd26, 8'd114}: color_data = 12'h249;
			{8'd26, 8'd115}: color_data = 12'h249;
			{8'd26, 8'd116}: color_data = 12'h249;
			{8'd26, 8'd117}: color_data = 12'h249;
			{8'd26, 8'd118}: color_data = 12'h249;
			{8'd26, 8'd119}: color_data = 12'h249;
			{8'd26, 8'd120}: color_data = 12'h249;
			{8'd26, 8'd121}: color_data = 12'h249;
			{8'd26, 8'd122}: color_data = 12'h249;
			{8'd26, 8'd123}: color_data = 12'h249;
			{8'd26, 8'd124}: color_data = 12'h249;
			{8'd26, 8'd125}: color_data = 12'h249;
			{8'd26, 8'd126}: color_data = 12'h249;
			{8'd26, 8'd127}: color_data = 12'h249;
			{8'd26, 8'd128}: color_data = 12'h249;
			{8'd26, 8'd129}: color_data = 12'h249;
			{8'd26, 8'd130}: color_data = 12'h249;
			{8'd26, 8'd131}: color_data = 12'h249;
			{8'd26, 8'd132}: color_data = 12'h249;
			{8'd26, 8'd133}: color_data = 12'h249;
			{8'd26, 8'd134}: color_data = 12'h249;
			{8'd26, 8'd135}: color_data = 12'h249;
			{8'd26, 8'd136}: color_data = 12'h249;
			{8'd26, 8'd137}: color_data = 12'h249;
			{8'd26, 8'd138}: color_data = 12'h224;
			{8'd26, 8'd139}: color_data = 12'h633;
			{8'd26, 8'd140}: color_data = 12'h633;
			{8'd26, 8'd141}: color_data = 12'h633;
			{8'd26, 8'd142}: color_data = 12'h643;
			{8'd26, 8'd143}: color_data = 12'h533;
			{8'd26, 8'd144}: color_data = 12'h643;
			{8'd26, 8'd145}: color_data = 12'h321;
			{8'd27, 8'd19}: color_data = 12'hfc5;
			{8'd27, 8'd20}: color_data = 12'hfc5;
			{8'd27, 8'd21}: color_data = 12'hfc4;
			{8'd27, 8'd22}: color_data = 12'hea1;
			{8'd27, 8'd23}: color_data = 12'heb3;
			{8'd27, 8'd24}: color_data = 12'hfc5;
			{8'd27, 8'd25}: color_data = 12'hfc6;
			{8'd27, 8'd26}: color_data = 12'hfc5;
			{8'd27, 8'd27}: color_data = 12'hfc5;
			{8'd27, 8'd28}: color_data = 12'hfc4;
			{8'd27, 8'd29}: color_data = 12'hfc5;
			{8'd27, 8'd30}: color_data = 12'hfc6;
			{8'd27, 8'd31}: color_data = 12'heb2;
			{8'd27, 8'd32}: color_data = 12'hd90;
			{8'd27, 8'd33}: color_data = 12'hd90;
			{8'd27, 8'd34}: color_data = 12'hd90;
			{8'd27, 8'd35}: color_data = 12'hfc4;
			{8'd27, 8'd36}: color_data = 12'hfc5;
			{8'd27, 8'd37}: color_data = 12'hfc5;
			{8'd27, 8'd50}: color_data = 12'h000;
			{8'd27, 8'd51}: color_data = 12'h062;
			{8'd27, 8'd52}: color_data = 12'h0a4;
			{8'd27, 8'd53}: color_data = 12'h0a3;
			{8'd27, 8'd54}: color_data = 12'h0a3;
			{8'd27, 8'd55}: color_data = 12'h0a3;
			{8'd27, 8'd56}: color_data = 12'h0a3;
			{8'd27, 8'd57}: color_data = 12'h0a3;
			{8'd27, 8'd58}: color_data = 12'h0a3;
			{8'd27, 8'd59}: color_data = 12'h0a3;
			{8'd27, 8'd60}: color_data = 12'h0a3;
			{8'd27, 8'd61}: color_data = 12'h0a3;
			{8'd27, 8'd62}: color_data = 12'h0a3;
			{8'd27, 8'd63}: color_data = 12'h093;
			{8'd27, 8'd64}: color_data = 12'h093;
			{8'd27, 8'd65}: color_data = 12'h093;
			{8'd27, 8'd66}: color_data = 12'h0a3;
			{8'd27, 8'd67}: color_data = 12'h0a3;
			{8'd27, 8'd68}: color_data = 12'h0a3;
			{8'd27, 8'd69}: color_data = 12'h093;
			{8'd27, 8'd70}: color_data = 12'h062;
			{8'd27, 8'd71}: color_data = 12'h0a3;
			{8'd27, 8'd72}: color_data = 12'h083;
			{8'd27, 8'd73}: color_data = 12'h987;
			{8'd27, 8'd74}: color_data = 12'hfdb;
			{8'd27, 8'd75}: color_data = 12'hfdb;
			{8'd27, 8'd76}: color_data = 12'hfdb;
			{8'd27, 8'd77}: color_data = 12'hfeb;
			{8'd27, 8'd78}: color_data = 12'h976;
			{8'd27, 8'd79}: color_data = 12'h521;
			{8'd27, 8'd80}: color_data = 12'h765;
			{8'd27, 8'd81}: color_data = 12'h754;
			{8'd27, 8'd82}: color_data = 12'ha87;
			{8'd27, 8'd83}: color_data = 12'hfdb;
			{8'd27, 8'd84}: color_data = 12'hfdb;
			{8'd27, 8'd85}: color_data = 12'hfdb;
			{8'd27, 8'd86}: color_data = 12'hfdb;
			{8'd27, 8'd87}: color_data = 12'h976;
			{8'd27, 8'd88}: color_data = 12'h742;
			{8'd27, 8'd89}: color_data = 12'h631;
			{8'd27, 8'd90}: color_data = 12'h000;
			{8'd27, 8'd91}: color_data = 12'h000;
			{8'd27, 8'd92}: color_data = 12'h124;
			{8'd27, 8'd93}: color_data = 12'h249;
			{8'd27, 8'd94}: color_data = 12'h249;
			{8'd27, 8'd95}: color_data = 12'h248;
			{8'd27, 8'd96}: color_data = 12'h345;
			{8'd27, 8'd97}: color_data = 12'h898;
			{8'd27, 8'd98}: color_data = 12'h133;
			{8'd27, 8'd99}: color_data = 12'h253;
			{8'd27, 8'd100}: color_data = 12'h797;
			{8'd27, 8'd101}: color_data = 12'h687;
			{8'd27, 8'd102}: color_data = 12'h173;
			{8'd27, 8'd103}: color_data = 12'h052;
			{8'd27, 8'd104}: color_data = 12'h136;
			{8'd27, 8'd105}: color_data = 12'h249;
			{8'd27, 8'd106}: color_data = 12'h249;
			{8'd27, 8'd107}: color_data = 12'h249;
			{8'd27, 8'd108}: color_data = 12'h249;
			{8'd27, 8'd109}: color_data = 12'h249;
			{8'd27, 8'd110}: color_data = 12'h249;
			{8'd27, 8'd111}: color_data = 12'h249;
			{8'd27, 8'd112}: color_data = 12'h249;
			{8'd27, 8'd113}: color_data = 12'h249;
			{8'd27, 8'd114}: color_data = 12'h249;
			{8'd27, 8'd115}: color_data = 12'h249;
			{8'd27, 8'd116}: color_data = 12'h249;
			{8'd27, 8'd117}: color_data = 12'h249;
			{8'd27, 8'd118}: color_data = 12'h249;
			{8'd27, 8'd119}: color_data = 12'h249;
			{8'd27, 8'd120}: color_data = 12'h249;
			{8'd27, 8'd121}: color_data = 12'h249;
			{8'd27, 8'd122}: color_data = 12'h249;
			{8'd27, 8'd123}: color_data = 12'h249;
			{8'd27, 8'd124}: color_data = 12'h249;
			{8'd27, 8'd125}: color_data = 12'h249;
			{8'd27, 8'd126}: color_data = 12'h249;
			{8'd27, 8'd127}: color_data = 12'h249;
			{8'd27, 8'd128}: color_data = 12'h249;
			{8'd27, 8'd129}: color_data = 12'h248;
			{8'd27, 8'd130}: color_data = 12'h136;
			{8'd27, 8'd131}: color_data = 12'h137;
			{8'd27, 8'd132}: color_data = 12'h249;
			{8'd27, 8'd133}: color_data = 12'h249;
			{8'd27, 8'd134}: color_data = 12'h249;
			{8'd27, 8'd135}: color_data = 12'h249;
			{8'd27, 8'd136}: color_data = 12'h249;
			{8'd27, 8'd137}: color_data = 12'h249;
			{8'd27, 8'd138}: color_data = 12'h224;
			{8'd27, 8'd139}: color_data = 12'h633;
			{8'd27, 8'd140}: color_data = 12'h633;
			{8'd27, 8'd141}: color_data = 12'h633;
			{8'd27, 8'd142}: color_data = 12'h633;
			{8'd27, 8'd143}: color_data = 12'h532;
			{8'd27, 8'd144}: color_data = 12'h432;
			{8'd28, 8'd19}: color_data = 12'hfc5;
			{8'd28, 8'd20}: color_data = 12'hfc5;
			{8'd28, 8'd21}: color_data = 12'heb2;
			{8'd28, 8'd22}: color_data = 12'hd90;
			{8'd28, 8'd23}: color_data = 12'hd90;
			{8'd28, 8'd24}: color_data = 12'hd90;
			{8'd28, 8'd25}: color_data = 12'hea0;
			{8'd28, 8'd26}: color_data = 12'heb2;
			{8'd28, 8'd27}: color_data = 12'hfb3;
			{8'd28, 8'd28}: color_data = 12'hfc5;
			{8'd28, 8'd29}: color_data = 12'hfc5;
			{8'd28, 8'd30}: color_data = 12'hfc6;
			{8'd28, 8'd31}: color_data = 12'hfc5;
			{8'd28, 8'd32}: color_data = 12'heb2;
			{8'd28, 8'd33}: color_data = 12'hd90;
			{8'd28, 8'd34}: color_data = 12'hda0;
			{8'd28, 8'd35}: color_data = 12'hfc5;
			{8'd28, 8'd36}: color_data = 12'hfc5;
			{8'd28, 8'd37}: color_data = 12'hfc5;
			{8'd28, 8'd50}: color_data = 12'h000;
			{8'd28, 8'd51}: color_data = 12'h072;
			{8'd28, 8'd52}: color_data = 12'h0a3;
			{8'd28, 8'd53}: color_data = 12'h0a3;
			{8'd28, 8'd54}: color_data = 12'h0a3;
			{8'd28, 8'd55}: color_data = 12'h0a3;
			{8'd28, 8'd56}: color_data = 12'h0a3;
			{8'd28, 8'd57}: color_data = 12'h0a3;
			{8'd28, 8'd58}: color_data = 12'h0a3;
			{8'd28, 8'd59}: color_data = 12'h0a3;
			{8'd28, 8'd60}: color_data = 12'h0a3;
			{8'd28, 8'd61}: color_data = 12'h093;
			{8'd28, 8'd62}: color_data = 12'h274;
			{8'd28, 8'd63}: color_data = 12'h797;
			{8'd28, 8'd64}: color_data = 12'h9a9;
			{8'd28, 8'd65}: color_data = 12'h898;
			{8'd28, 8'd66}: color_data = 12'h375;
			{8'd28, 8'd67}: color_data = 12'h093;
			{8'd28, 8'd68}: color_data = 12'h083;
			{8'd28, 8'd69}: color_data = 12'h062;
			{8'd28, 8'd70}: color_data = 12'h0a3;
			{8'd28, 8'd71}: color_data = 12'h0a3;
			{8'd28, 8'd72}: color_data = 12'h163;
			{8'd28, 8'd73}: color_data = 12'ha87;
			{8'd28, 8'd74}: color_data = 12'ha97;
			{8'd28, 8'd75}: color_data = 12'ha97;
			{8'd28, 8'd76}: color_data = 12'hfdb;
			{8'd28, 8'd77}: color_data = 12'hfdb;
			{8'd28, 8'd78}: color_data = 12'hca9;
			{8'd28, 8'd79}: color_data = 12'ha87;
			{8'd28, 8'd80}: color_data = 12'hfdb;
			{8'd28, 8'd81}: color_data = 12'hfdb;
			{8'd28, 8'd82}: color_data = 12'hfdb;
			{8'd28, 8'd83}: color_data = 12'hfdb;
			{8'd28, 8'd84}: color_data = 12'hfdb;
			{8'd28, 8'd85}: color_data = 12'hfdb;
			{8'd28, 8'd86}: color_data = 12'hfdb;
			{8'd28, 8'd87}: color_data = 12'heca;
			{8'd28, 8'd88}: color_data = 12'h432;
			{8'd28, 8'd89}: color_data = 12'h100;
			{8'd28, 8'd91}: color_data = 12'h013;
			{8'd28, 8'd92}: color_data = 12'h249;
			{8'd28, 8'd93}: color_data = 12'h249;
			{8'd28, 8'd94}: color_data = 12'h136;
			{8'd28, 8'd95}: color_data = 12'h053;
			{8'd28, 8'd96}: color_data = 12'h083;
			{8'd28, 8'd97}: color_data = 12'h092;
			{8'd28, 8'd98}: color_data = 12'h0a3;
			{8'd28, 8'd99}: color_data = 12'h0a3;
			{8'd28, 8'd100}: color_data = 12'h093;
			{8'd28, 8'd101}: color_data = 12'h093;
			{8'd28, 8'd102}: color_data = 12'h0a3;
			{8'd28, 8'd103}: color_data = 12'h053;
			{8'd28, 8'd104}: color_data = 12'h249;
			{8'd28, 8'd105}: color_data = 12'h249;
			{8'd28, 8'd106}: color_data = 12'h249;
			{8'd28, 8'd107}: color_data = 12'h249;
			{8'd28, 8'd108}: color_data = 12'h249;
			{8'd28, 8'd109}: color_data = 12'h249;
			{8'd28, 8'd110}: color_data = 12'h249;
			{8'd28, 8'd111}: color_data = 12'h249;
			{8'd28, 8'd112}: color_data = 12'h249;
			{8'd28, 8'd113}: color_data = 12'h249;
			{8'd28, 8'd114}: color_data = 12'h249;
			{8'd28, 8'd115}: color_data = 12'h249;
			{8'd28, 8'd116}: color_data = 12'h249;
			{8'd28, 8'd117}: color_data = 12'h249;
			{8'd28, 8'd118}: color_data = 12'h249;
			{8'd28, 8'd119}: color_data = 12'h249;
			{8'd28, 8'd120}: color_data = 12'h249;
			{8'd28, 8'd121}: color_data = 12'h249;
			{8'd28, 8'd122}: color_data = 12'h249;
			{8'd28, 8'd123}: color_data = 12'h249;
			{8'd28, 8'd124}: color_data = 12'h249;
			{8'd28, 8'd125}: color_data = 12'h249;
			{8'd28, 8'd126}: color_data = 12'h248;
			{8'd28, 8'd127}: color_data = 12'h136;
			{8'd28, 8'd128}: color_data = 12'h124;
			{8'd28, 8'd129}: color_data = 12'h012;
			{8'd28, 8'd130}: color_data = 12'h000;
			{8'd28, 8'd131}: color_data = 12'h124;
			{8'd28, 8'd132}: color_data = 12'h136;
			{8'd28, 8'd133}: color_data = 12'h249;
			{8'd28, 8'd134}: color_data = 12'h249;
			{8'd28, 8'd135}: color_data = 12'h249;
			{8'd28, 8'd136}: color_data = 12'h249;
			{8'd28, 8'd137}: color_data = 12'h249;
			{8'd28, 8'd138}: color_data = 12'h223;
			{8'd28, 8'd139}: color_data = 12'h633;
			{8'd28, 8'd140}: color_data = 12'h633;
			{8'd28, 8'd141}: color_data = 12'h633;
			{8'd28, 8'd142}: color_data = 12'h633;
			{8'd28, 8'd143}: color_data = 12'h532;
			{8'd28, 8'd144}: color_data = 12'h221;
			{8'd29, 8'd18}: color_data = 12'hfd6;
			{8'd29, 8'd19}: color_data = 12'hfc5;
			{8'd29, 8'd20}: color_data = 12'hfc5;
			{8'd29, 8'd21}: color_data = 12'hea0;
			{8'd29, 8'd22}: color_data = 12'hd90;
			{8'd29, 8'd23}: color_data = 12'hd90;
			{8'd29, 8'd24}: color_data = 12'hd90;
			{8'd29, 8'd25}: color_data = 12'hd90;
			{8'd29, 8'd26}: color_data = 12'hd90;
			{8'd29, 8'd27}: color_data = 12'hd90;
			{8'd29, 8'd28}: color_data = 12'hda0;
			{8'd29, 8'd29}: color_data = 12'hea1;
			{8'd29, 8'd30}: color_data = 12'heb3;
			{8'd29, 8'd31}: color_data = 12'hfc5;
			{8'd29, 8'd32}: color_data = 12'hfc5;
			{8'd29, 8'd33}: color_data = 12'heb2;
			{8'd29, 8'd34}: color_data = 12'heb1;
			{8'd29, 8'd35}: color_data = 12'hfc5;
			{8'd29, 8'd36}: color_data = 12'hfc5;
			{8'd29, 8'd37}: color_data = 12'hfa5;
			{8'd29, 8'd50}: color_data = 12'h000;
			{8'd29, 8'd51}: color_data = 12'h072;
			{8'd29, 8'd52}: color_data = 12'h0a3;
			{8'd29, 8'd53}: color_data = 12'h0a3;
			{8'd29, 8'd54}: color_data = 12'h0a3;
			{8'd29, 8'd55}: color_data = 12'h0a3;
			{8'd29, 8'd56}: color_data = 12'h0a3;
			{8'd29, 8'd57}: color_data = 12'h0a3;
			{8'd29, 8'd58}: color_data = 12'h0a3;
			{8'd29, 8'd59}: color_data = 12'h0a3;
			{8'd29, 8'd60}: color_data = 12'h083;
			{8'd29, 8'd61}: color_data = 12'h787;
			{8'd29, 8'd62}: color_data = 12'hfee;
			{8'd29, 8'd63}: color_data = 12'hfff;
			{8'd29, 8'd64}: color_data = 12'hfff;
			{8'd29, 8'd65}: color_data = 12'hfff;
			{8'd29, 8'd66}: color_data = 12'hfff;
			{8'd29, 8'd67}: color_data = 12'h676;
			{8'd29, 8'd68}: color_data = 12'h051;
			{8'd29, 8'd69}: color_data = 12'h0a3;
			{8'd29, 8'd70}: color_data = 12'h0a3;
			{8'd29, 8'd71}: color_data = 12'h082;
			{8'd29, 8'd72}: color_data = 12'h665;
			{8'd29, 8'd73}: color_data = 12'hdb9;
			{8'd29, 8'd74}: color_data = 12'heca;
			{8'd29, 8'd75}: color_data = 12'hfdb;
			{8'd29, 8'd76}: color_data = 12'hfdb;
			{8'd29, 8'd77}: color_data = 12'hfdb;
			{8'd29, 8'd78}: color_data = 12'hfdb;
			{8'd29, 8'd79}: color_data = 12'hfeb;
			{8'd29, 8'd80}: color_data = 12'hfdb;
			{8'd29, 8'd81}: color_data = 12'hfdb;
			{8'd29, 8'd82}: color_data = 12'hfdb;
			{8'd29, 8'd83}: color_data = 12'hfdb;
			{8'd29, 8'd84}: color_data = 12'hfdb;
			{8'd29, 8'd85}: color_data = 12'hfdb;
			{8'd29, 8'd86}: color_data = 12'hfdb;
			{8'd29, 8'd87}: color_data = 12'hfeb;
			{8'd29, 8'd88}: color_data = 12'h987;
			{8'd29, 8'd89}: color_data = 12'h000;
			{8'd29, 8'd90}: color_data = 12'h001;
			{8'd29, 8'd91}: color_data = 12'h248;
			{8'd29, 8'd92}: color_data = 12'h249;
			{8'd29, 8'd93}: color_data = 12'h044;
			{8'd29, 8'd94}: color_data = 12'h082;
			{8'd29, 8'd95}: color_data = 12'h0a3;
			{8'd29, 8'd96}: color_data = 12'h0a3;
			{8'd29, 8'd97}: color_data = 12'h0a3;
			{8'd29, 8'd98}: color_data = 12'h0a3;
			{8'd29, 8'd99}: color_data = 12'h0a3;
			{8'd29, 8'd100}: color_data = 12'h0a3;
			{8'd29, 8'd101}: color_data = 12'h0a3;
			{8'd29, 8'd102}: color_data = 12'h0a3;
			{8'd29, 8'd103}: color_data = 12'h145;
			{8'd29, 8'd104}: color_data = 12'h249;
			{8'd29, 8'd105}: color_data = 12'h249;
			{8'd29, 8'd106}: color_data = 12'h249;
			{8'd29, 8'd107}: color_data = 12'h249;
			{8'd29, 8'd108}: color_data = 12'h249;
			{8'd29, 8'd109}: color_data = 12'h249;
			{8'd29, 8'd110}: color_data = 12'h249;
			{8'd29, 8'd111}: color_data = 12'h249;
			{8'd29, 8'd112}: color_data = 12'h249;
			{8'd29, 8'd113}: color_data = 12'h249;
			{8'd29, 8'd114}: color_data = 12'h249;
			{8'd29, 8'd115}: color_data = 12'h249;
			{8'd29, 8'd116}: color_data = 12'h249;
			{8'd29, 8'd117}: color_data = 12'h249;
			{8'd29, 8'd118}: color_data = 12'h249;
			{8'd29, 8'd119}: color_data = 12'h249;
			{8'd29, 8'd120}: color_data = 12'h249;
			{8'd29, 8'd121}: color_data = 12'h249;
			{8'd29, 8'd122}: color_data = 12'h249;
			{8'd29, 8'd123}: color_data = 12'h249;
			{8'd29, 8'd124}: color_data = 12'h249;
			{8'd29, 8'd125}: color_data = 12'h136;
			{8'd29, 8'd126}: color_data = 12'h012;
			{8'd29, 8'd127}: color_data = 12'h000;
			{8'd29, 8'd131}: color_data = 12'h000;
			{8'd29, 8'd132}: color_data = 12'h001;
			{8'd29, 8'd133}: color_data = 12'h247;
			{8'd29, 8'd134}: color_data = 12'h249;
			{8'd29, 8'd135}: color_data = 12'h249;
			{8'd29, 8'd136}: color_data = 12'h249;
			{8'd29, 8'd137}: color_data = 12'h249;
			{8'd29, 8'd138}: color_data = 12'h323;
			{8'd29, 8'd139}: color_data = 12'h643;
			{8'd29, 8'd140}: color_data = 12'h633;
			{8'd29, 8'd141}: color_data = 12'h643;
			{8'd29, 8'd142}: color_data = 12'h533;
			{8'd29, 8'd143}: color_data = 12'h432;
			{8'd29, 8'd144}: color_data = 12'h000;
			{8'd30, 8'd18}: color_data = 12'hfc6;
			{8'd30, 8'd19}: color_data = 12'hfc5;
			{8'd30, 8'd20}: color_data = 12'hfc4;
			{8'd30, 8'd21}: color_data = 12'hd90;
			{8'd30, 8'd22}: color_data = 12'hd90;
			{8'd30, 8'd23}: color_data = 12'hd90;
			{8'd30, 8'd24}: color_data = 12'hd90;
			{8'd30, 8'd25}: color_data = 12'hd90;
			{8'd30, 8'd26}: color_data = 12'hd90;
			{8'd30, 8'd27}: color_data = 12'hd90;
			{8'd30, 8'd28}: color_data = 12'hd90;
			{8'd30, 8'd29}: color_data = 12'hd90;
			{8'd30, 8'd30}: color_data = 12'hd90;
			{8'd30, 8'd31}: color_data = 12'hd90;
			{8'd30, 8'd32}: color_data = 12'hea1;
			{8'd30, 8'd33}: color_data = 12'heb2;
			{8'd30, 8'd34}: color_data = 12'hfc4;
			{8'd30, 8'd35}: color_data = 12'hfc5;
			{8'd30, 8'd36}: color_data = 12'hfc4;
			{8'd30, 8'd50}: color_data = 12'h000;
			{8'd30, 8'd51}: color_data = 12'h062;
			{8'd30, 8'd52}: color_data = 12'h0a4;
			{8'd30, 8'd53}: color_data = 12'h0a3;
			{8'd30, 8'd54}: color_data = 12'h0a3;
			{8'd30, 8'd55}: color_data = 12'h0a3;
			{8'd30, 8'd56}: color_data = 12'h0a3;
			{8'd30, 8'd57}: color_data = 12'h0a3;
			{8'd30, 8'd58}: color_data = 12'h0a3;
			{8'd30, 8'd59}: color_data = 12'h0a3;
			{8'd30, 8'd60}: color_data = 12'h586;
			{8'd30, 8'd61}: color_data = 12'hfff;
			{8'd30, 8'd62}: color_data = 12'hefe;
			{8'd30, 8'd63}: color_data = 12'hefe;
			{8'd30, 8'd64}: color_data = 12'hfff;
			{8'd30, 8'd65}: color_data = 12'hfff;
			{8'd30, 8'd66}: color_data = 12'heee;
			{8'd30, 8'd67}: color_data = 12'h375;
			{8'd30, 8'd68}: color_data = 12'h0a3;
			{8'd30, 8'd69}: color_data = 12'h0a3;
			{8'd30, 8'd70}: color_data = 12'h0a3;
			{8'd30, 8'd71}: color_data = 12'h363;
			{8'd30, 8'd72}: color_data = 12'hca8;
			{8'd30, 8'd73}: color_data = 12'hca8;
			{8'd30, 8'd74}: color_data = 12'ha97;
			{8'd30, 8'd75}: color_data = 12'h987;
			{8'd30, 8'd76}: color_data = 12'ha97;
			{8'd30, 8'd77}: color_data = 12'hfdb;
			{8'd30, 8'd78}: color_data = 12'hfdb;
			{8'd30, 8'd79}: color_data = 12'hfdb;
			{8'd30, 8'd80}: color_data = 12'hfdb;
			{8'd30, 8'd81}: color_data = 12'h987;
			{8'd30, 8'd82}: color_data = 12'hba8;
			{8'd30, 8'd83}: color_data = 12'hfdb;
			{8'd30, 8'd84}: color_data = 12'hfdb;
			{8'd30, 8'd85}: color_data = 12'hfdb;
			{8'd30, 8'd86}: color_data = 12'hfdb;
			{8'd30, 8'd87}: color_data = 12'hfdb;
			{8'd30, 8'd88}: color_data = 12'hdb9;
			{8'd30, 8'd89}: color_data = 12'h100;
			{8'd30, 8'd90}: color_data = 12'h125;
			{8'd30, 8'd91}: color_data = 12'h249;
			{8'd30, 8'd92}: color_data = 12'h034;
			{8'd30, 8'd93}: color_data = 12'h093;
			{8'd30, 8'd94}: color_data = 12'h0a3;
			{8'd30, 8'd95}: color_data = 12'h0a3;
			{8'd30, 8'd96}: color_data = 12'h0a3;
			{8'd30, 8'd97}: color_data = 12'h0a3;
			{8'd30, 8'd98}: color_data = 12'h0a3;
			{8'd30, 8'd99}: color_data = 12'h0a3;
			{8'd30, 8'd100}: color_data = 12'h0a3;
			{8'd30, 8'd101}: color_data = 12'h0a3;
			{8'd30, 8'd102}: color_data = 12'h093;
			{8'd30, 8'd103}: color_data = 12'h136;
			{8'd30, 8'd104}: color_data = 12'h249;
			{8'd30, 8'd105}: color_data = 12'h249;
			{8'd30, 8'd106}: color_data = 12'h249;
			{8'd30, 8'd107}: color_data = 12'h249;
			{8'd30, 8'd108}: color_data = 12'h249;
			{8'd30, 8'd109}: color_data = 12'h249;
			{8'd30, 8'd110}: color_data = 12'h249;
			{8'd30, 8'd111}: color_data = 12'h249;
			{8'd30, 8'd112}: color_data = 12'h249;
			{8'd30, 8'd113}: color_data = 12'h249;
			{8'd30, 8'd114}: color_data = 12'h249;
			{8'd30, 8'd115}: color_data = 12'h249;
			{8'd30, 8'd116}: color_data = 12'h249;
			{8'd30, 8'd117}: color_data = 12'h249;
			{8'd30, 8'd118}: color_data = 12'h249;
			{8'd30, 8'd119}: color_data = 12'h249;
			{8'd30, 8'd120}: color_data = 12'h249;
			{8'd30, 8'd121}: color_data = 12'h249;
			{8'd30, 8'd122}: color_data = 12'h249;
			{8'd30, 8'd123}: color_data = 12'h248;
			{8'd30, 8'd124}: color_data = 12'h013;
			{8'd30, 8'd125}: color_data = 12'h000;
			{8'd30, 8'd133}: color_data = 12'h013;
			{8'd30, 8'd134}: color_data = 12'h248;
			{8'd30, 8'd135}: color_data = 12'h249;
			{8'd30, 8'd136}: color_data = 12'h249;
			{8'd30, 8'd137}: color_data = 12'h147;
			{8'd30, 8'd138}: color_data = 12'h422;
			{8'd30, 8'd139}: color_data = 12'h643;
			{8'd30, 8'd140}: color_data = 12'h633;
			{8'd30, 8'd141}: color_data = 12'h643;
			{8'd30, 8'd142}: color_data = 12'h533;
			{8'd30, 8'd143}: color_data = 12'h331;
			{8'd30, 8'd144}: color_data = 12'h000;
			{8'd31, 8'd18}: color_data = 12'hfc5;
			{8'd31, 8'd19}: color_data = 12'hfc5;
			{8'd31, 8'd20}: color_data = 12'heb3;
			{8'd31, 8'd21}: color_data = 12'hd90;
			{8'd31, 8'd22}: color_data = 12'hd90;
			{8'd31, 8'd23}: color_data = 12'hd90;
			{8'd31, 8'd24}: color_data = 12'hd90;
			{8'd31, 8'd25}: color_data = 12'hd90;
			{8'd31, 8'd26}: color_data = 12'hd90;
			{8'd31, 8'd27}: color_data = 12'hd90;
			{8'd31, 8'd28}: color_data = 12'hd90;
			{8'd31, 8'd29}: color_data = 12'hd90;
			{8'd31, 8'd30}: color_data = 12'hd90;
			{8'd31, 8'd31}: color_data = 12'hd90;
			{8'd31, 8'd32}: color_data = 12'hd90;
			{8'd31, 8'd33}: color_data = 12'hd90;
			{8'd31, 8'd34}: color_data = 12'hfb3;
			{8'd31, 8'd35}: color_data = 12'hfc5;
			{8'd31, 8'd36}: color_data = 12'hfc4;
			{8'd31, 8'd51}: color_data = 12'h031;
			{8'd31, 8'd52}: color_data = 12'h093;
			{8'd31, 8'd53}: color_data = 12'h0a3;
			{8'd31, 8'd54}: color_data = 12'h0a3;
			{8'd31, 8'd55}: color_data = 12'h0a3;
			{8'd31, 8'd56}: color_data = 12'h0a3;
			{8'd31, 8'd57}: color_data = 12'h0a3;
			{8'd31, 8'd58}: color_data = 12'h0a3;
			{8'd31, 8'd59}: color_data = 12'h092;
			{8'd31, 8'd60}: color_data = 12'h9aa;
			{8'd31, 8'd61}: color_data = 12'hfff;
			{8'd31, 8'd62}: color_data = 12'hced;
			{8'd31, 8'd63}: color_data = 12'haeb;
			{8'd31, 8'd64}: color_data = 12'h9eb;
			{8'd31, 8'd65}: color_data = 12'h9ca;
			{8'd31, 8'd66}: color_data = 12'h475;
			{8'd31, 8'd67}: color_data = 12'h093;
			{8'd31, 8'd68}: color_data = 12'h0a3;
			{8'd31, 8'd69}: color_data = 12'h0a3;
			{8'd31, 8'd70}: color_data = 12'h072;
			{8'd31, 8'd71}: color_data = 12'h876;
			{8'd31, 8'd72}: color_data = 12'hfec;
			{8'd31, 8'd73}: color_data = 12'hfdb;
			{8'd31, 8'd74}: color_data = 12'hfdb;
			{8'd31, 8'd75}: color_data = 12'hfdb;
			{8'd31, 8'd76}: color_data = 12'hba8;
			{8'd31, 8'd77}: color_data = 12'h765;
			{8'd31, 8'd78}: color_data = 12'hdca;
			{8'd31, 8'd79}: color_data = 12'hfdb;
			{8'd31, 8'd80}: color_data = 12'hfeb;
			{8'd31, 8'd81}: color_data = 12'h765;
			{8'd31, 8'd82}: color_data = 12'h110;
			{8'd31, 8'd83}: color_data = 12'heca;
			{8'd31, 8'd84}: color_data = 12'hfdb;
			{8'd31, 8'd85}: color_data = 12'hfdb;
			{8'd31, 8'd86}: color_data = 12'hfdb;
			{8'd31, 8'd87}: color_data = 12'hfdb;
			{8'd31, 8'd88}: color_data = 12'hfdb;
			{8'd31, 8'd89}: color_data = 12'h322;
			{8'd31, 8'd90}: color_data = 12'h036;
			{8'd31, 8'd91}: color_data = 12'h346;
			{8'd31, 8'd92}: color_data = 12'h464;
			{8'd31, 8'd93}: color_data = 12'h0a3;
			{8'd31, 8'd94}: color_data = 12'h0a3;
			{8'd31, 8'd95}: color_data = 12'h0a3;
			{8'd31, 8'd96}: color_data = 12'h0a3;
			{8'd31, 8'd97}: color_data = 12'h0a3;
			{8'd31, 8'd98}: color_data = 12'h0a3;
			{8'd31, 8'd99}: color_data = 12'h0a3;
			{8'd31, 8'd100}: color_data = 12'h0a3;
			{8'd31, 8'd101}: color_data = 12'h0a3;
			{8'd31, 8'd102}: color_data = 12'h083;
			{8'd31, 8'd103}: color_data = 12'h137;
			{8'd31, 8'd104}: color_data = 12'h249;
			{8'd31, 8'd105}: color_data = 12'h249;
			{8'd31, 8'd106}: color_data = 12'h249;
			{8'd31, 8'd107}: color_data = 12'h249;
			{8'd31, 8'd108}: color_data = 12'h249;
			{8'd31, 8'd109}: color_data = 12'h249;
			{8'd31, 8'd110}: color_data = 12'h249;
			{8'd31, 8'd111}: color_data = 12'h249;
			{8'd31, 8'd112}: color_data = 12'h249;
			{8'd31, 8'd113}: color_data = 12'h249;
			{8'd31, 8'd114}: color_data = 12'h249;
			{8'd31, 8'd115}: color_data = 12'h249;
			{8'd31, 8'd116}: color_data = 12'h249;
			{8'd31, 8'd117}: color_data = 12'h249;
			{8'd31, 8'd118}: color_data = 12'h249;
			{8'd31, 8'd119}: color_data = 12'h249;
			{8'd31, 8'd120}: color_data = 12'h249;
			{8'd31, 8'd121}: color_data = 12'h249;
			{8'd31, 8'd122}: color_data = 12'h249;
			{8'd31, 8'd123}: color_data = 12'h125;
			{8'd31, 8'd124}: color_data = 12'h000;
			{8'd31, 8'd133}: color_data = 12'h000;
			{8'd31, 8'd134}: color_data = 12'h124;
			{8'd31, 8'd135}: color_data = 12'h248;
			{8'd31, 8'd136}: color_data = 12'h249;
			{8'd31, 8'd137}: color_data = 12'h224;
			{8'd31, 8'd138}: color_data = 12'h633;
			{8'd31, 8'd139}: color_data = 12'h633;
			{8'd31, 8'd140}: color_data = 12'h633;
			{8'd31, 8'd141}: color_data = 12'h643;
			{8'd31, 8'd142}: color_data = 12'h432;
			{8'd31, 8'd143}: color_data = 12'h321;
			{8'd32, 8'd17}: color_data = 12'hfff;
			{8'd32, 8'd18}: color_data = 12'hfc4;
			{8'd32, 8'd19}: color_data = 12'hfc5;
			{8'd32, 8'd20}: color_data = 12'hea1;
			{8'd32, 8'd21}: color_data = 12'hd90;
			{8'd32, 8'd22}: color_data = 12'hd90;
			{8'd32, 8'd23}: color_data = 12'hd90;
			{8'd32, 8'd24}: color_data = 12'heb2;
			{8'd32, 8'd25}: color_data = 12'heb2;
			{8'd32, 8'd26}: color_data = 12'hea1;
			{8'd32, 8'd27}: color_data = 12'hd90;
			{8'd32, 8'd28}: color_data = 12'hd90;
			{8'd32, 8'd29}: color_data = 12'hd90;
			{8'd32, 8'd30}: color_data = 12'hd90;
			{8'd32, 8'd31}: color_data = 12'hd90;
			{8'd32, 8'd32}: color_data = 12'hd90;
			{8'd32, 8'd33}: color_data = 12'hd90;
			{8'd32, 8'd34}: color_data = 12'hfc4;
			{8'd32, 8'd35}: color_data = 12'hfc5;
			{8'd32, 8'd36}: color_data = 12'hfc5;
			{8'd32, 8'd51}: color_data = 12'h000;
			{8'd32, 8'd52}: color_data = 12'h041;
			{8'd32, 8'd53}: color_data = 12'h093;
			{8'd32, 8'd54}: color_data = 12'h0a3;
			{8'd32, 8'd55}: color_data = 12'h0a3;
			{8'd32, 8'd56}: color_data = 12'h0a3;
			{8'd32, 8'd57}: color_data = 12'h0a3;
			{8'd32, 8'd58}: color_data = 12'h0a3;
			{8'd32, 8'd59}: color_data = 12'h093;
			{8'd32, 8'd60}: color_data = 12'h797;
			{8'd32, 8'd61}: color_data = 12'hfff;
			{8'd32, 8'd62}: color_data = 12'hfff;
			{8'd32, 8'd63}: color_data = 12'hfff;
			{8'd32, 8'd64}: color_data = 12'h8ba;
			{8'd32, 8'd65}: color_data = 12'h163;
			{8'd32, 8'd66}: color_data = 12'h093;
			{8'd32, 8'd67}: color_data = 12'h0a3;
			{8'd32, 8'd68}: color_data = 12'h0a3;
			{8'd32, 8'd69}: color_data = 12'h093;
			{8'd32, 8'd70}: color_data = 12'h786;
			{8'd32, 8'd71}: color_data = 12'ha87;
			{8'd32, 8'd72}: color_data = 12'hfdb;
			{8'd32, 8'd73}: color_data = 12'hfdb;
			{8'd32, 8'd74}: color_data = 12'hfdb;
			{8'd32, 8'd75}: color_data = 12'ha97;
			{8'd32, 8'd76}: color_data = 12'h222;
			{8'd32, 8'd77}: color_data = 12'h876;
			{8'd32, 8'd78}: color_data = 12'heca;
			{8'd32, 8'd79}: color_data = 12'hfdb;
			{8'd32, 8'd80}: color_data = 12'hfeb;
			{8'd32, 8'd81}: color_data = 12'hba8;
			{8'd32, 8'd82}: color_data = 12'h000;
			{8'd32, 8'd83}: color_data = 12'ha97;
			{8'd32, 8'd84}: color_data = 12'hfeb;
			{8'd32, 8'd85}: color_data = 12'hfdb;
			{8'd32, 8'd86}: color_data = 12'hfdb;
			{8'd32, 8'd87}: color_data = 12'hfdb;
			{8'd32, 8'd88}: color_data = 12'hfdb;
			{8'd32, 8'd89}: color_data = 12'h765;
			{8'd32, 8'd90}: color_data = 12'h877;
			{8'd32, 8'd91}: color_data = 12'heca;
			{8'd32, 8'd92}: color_data = 12'hba8;
			{8'd32, 8'd93}: color_data = 12'h083;
			{8'd32, 8'd94}: color_data = 12'h0a3;
			{8'd32, 8'd95}: color_data = 12'h0a3;
			{8'd32, 8'd96}: color_data = 12'h0a3;
			{8'd32, 8'd97}: color_data = 12'h0a3;
			{8'd32, 8'd98}: color_data = 12'h0a3;
			{8'd32, 8'd99}: color_data = 12'h0a3;
			{8'd32, 8'd100}: color_data = 12'h0a3;
			{8'd32, 8'd101}: color_data = 12'h0a3;
			{8'd32, 8'd102}: color_data = 12'h073;
			{8'd32, 8'd103}: color_data = 12'h237;
			{8'd32, 8'd104}: color_data = 12'h249;
			{8'd32, 8'd105}: color_data = 12'h249;
			{8'd32, 8'd106}: color_data = 12'h249;
			{8'd32, 8'd107}: color_data = 12'h249;
			{8'd32, 8'd108}: color_data = 12'h249;
			{8'd32, 8'd109}: color_data = 12'h249;
			{8'd32, 8'd110}: color_data = 12'h249;
			{8'd32, 8'd111}: color_data = 12'h249;
			{8'd32, 8'd112}: color_data = 12'h249;
			{8'd32, 8'd113}: color_data = 12'h249;
			{8'd32, 8'd114}: color_data = 12'h249;
			{8'd32, 8'd115}: color_data = 12'h249;
			{8'd32, 8'd116}: color_data = 12'h249;
			{8'd32, 8'd117}: color_data = 12'h249;
			{8'd32, 8'd118}: color_data = 12'h249;
			{8'd32, 8'd119}: color_data = 12'h249;
			{8'd32, 8'd120}: color_data = 12'h249;
			{8'd32, 8'd121}: color_data = 12'h249;
			{8'd32, 8'd122}: color_data = 12'h248;
			{8'd32, 8'd123}: color_data = 12'h012;
			{8'd32, 8'd134}: color_data = 12'h000;
			{8'd32, 8'd135}: color_data = 12'h013;
			{8'd32, 8'd136}: color_data = 12'h123;
			{8'd32, 8'd137}: color_data = 12'h532;
			{8'd32, 8'd138}: color_data = 12'h643;
			{8'd32, 8'd139}: color_data = 12'h633;
			{8'd32, 8'd140}: color_data = 12'h643;
			{8'd32, 8'd141}: color_data = 12'h532;
			{8'd32, 8'd142}: color_data = 12'h100;
			{8'd32, 8'd143}: color_data = 12'h000;
			{8'd33, 8'd17}: color_data = 12'hfc5;
			{8'd33, 8'd18}: color_data = 12'hfc5;
			{8'd33, 8'd19}: color_data = 12'hfc4;
			{8'd33, 8'd20}: color_data = 12'hea0;
			{8'd33, 8'd21}: color_data = 12'hd90;
			{8'd33, 8'd22}: color_data = 12'hd90;
			{8'd33, 8'd23}: color_data = 12'hd90;
			{8'd33, 8'd24}: color_data = 12'hfb3;
			{8'd33, 8'd25}: color_data = 12'hfd7;
			{8'd33, 8'd26}: color_data = 12'hfb3;
			{8'd33, 8'd27}: color_data = 12'hd90;
			{8'd33, 8'd28}: color_data = 12'hd90;
			{8'd33, 8'd29}: color_data = 12'hd90;
			{8'd33, 8'd30}: color_data = 12'hda0;
			{8'd33, 8'd31}: color_data = 12'hea0;
			{8'd33, 8'd32}: color_data = 12'hd90;
			{8'd33, 8'd33}: color_data = 12'hd90;
			{8'd33, 8'd34}: color_data = 12'hfc4;
			{8'd33, 8'd35}: color_data = 12'hfc5;
			{8'd33, 8'd36}: color_data = 12'hfc5;
			{8'd33, 8'd52}: color_data = 12'h000;
			{8'd33, 8'd53}: color_data = 12'h020;
			{8'd33, 8'd54}: color_data = 12'h052;
			{8'd33, 8'd55}: color_data = 12'h072;
			{8'd33, 8'd56}: color_data = 12'h072;
			{8'd33, 8'd57}: color_data = 12'h083;
			{8'd33, 8'd58}: color_data = 12'h083;
			{8'd33, 8'd59}: color_data = 12'h083;
			{8'd33, 8'd60}: color_data = 12'h062;
			{8'd33, 8'd61}: color_data = 12'h454;
			{8'd33, 8'd62}: color_data = 12'h676;
			{8'd33, 8'd63}: color_data = 12'h697;
			{8'd33, 8'd64}: color_data = 12'h173;
			{8'd33, 8'd65}: color_data = 12'h0a3;
			{8'd33, 8'd66}: color_data = 12'h0a3;
			{8'd33, 8'd67}: color_data = 12'h0a3;
			{8'd33, 8'd68}: color_data = 12'h0a3;
			{8'd33, 8'd69}: color_data = 12'h252;
			{8'd33, 8'd70}: color_data = 12'h987;
			{8'd33, 8'd71}: color_data = 12'h876;
			{8'd33, 8'd72}: color_data = 12'h875;
			{8'd33, 8'd73}: color_data = 12'hfdb;
			{8'd33, 8'd74}: color_data = 12'hfdb;
			{8'd33, 8'd75}: color_data = 12'h433;
			{8'd33, 8'd76}: color_data = 12'hca9;
			{8'd33, 8'd77}: color_data = 12'hfec;
			{8'd33, 8'd78}: color_data = 12'hfdb;
			{8'd33, 8'd79}: color_data = 12'hfdb;
			{8'd33, 8'd80}: color_data = 12'hfdb;
			{8'd33, 8'd81}: color_data = 12'hcb9;
			{8'd33, 8'd82}: color_data = 12'h000;
			{8'd33, 8'd83}: color_data = 12'h654;
			{8'd33, 8'd84}: color_data = 12'hfdb;
			{8'd33, 8'd85}: color_data = 12'hfdb;
			{8'd33, 8'd86}: color_data = 12'hfdb;
			{8'd33, 8'd87}: color_data = 12'hfdb;
			{8'd33, 8'd88}: color_data = 12'hfdb;
			{8'd33, 8'd89}: color_data = 12'ha97;
			{8'd33, 8'd90}: color_data = 12'hfdb;
			{8'd33, 8'd91}: color_data = 12'hfeb;
			{8'd33, 8'd92}: color_data = 12'hca9;
			{8'd33, 8'd93}: color_data = 12'h083;
			{8'd33, 8'd94}: color_data = 12'h0a3;
			{8'd33, 8'd95}: color_data = 12'h0a3;
			{8'd33, 8'd96}: color_data = 12'h0a3;
			{8'd33, 8'd97}: color_data = 12'h0a3;
			{8'd33, 8'd98}: color_data = 12'h0a3;
			{8'd33, 8'd99}: color_data = 12'h0a3;
			{8'd33, 8'd100}: color_data = 12'h0a3;
			{8'd33, 8'd101}: color_data = 12'h0b3;
			{8'd33, 8'd102}: color_data = 12'h073;
			{8'd33, 8'd103}: color_data = 12'h238;
			{8'd33, 8'd104}: color_data = 12'h249;
			{8'd33, 8'd105}: color_data = 12'h249;
			{8'd33, 8'd106}: color_data = 12'h249;
			{8'd33, 8'd107}: color_data = 12'h249;
			{8'd33, 8'd108}: color_data = 12'h249;
			{8'd33, 8'd109}: color_data = 12'h249;
			{8'd33, 8'd110}: color_data = 12'h249;
			{8'd33, 8'd111}: color_data = 12'h249;
			{8'd33, 8'd112}: color_data = 12'h249;
			{8'd33, 8'd113}: color_data = 12'h249;
			{8'd33, 8'd114}: color_data = 12'h249;
			{8'd33, 8'd115}: color_data = 12'h249;
			{8'd33, 8'd116}: color_data = 12'h249;
			{8'd33, 8'd117}: color_data = 12'h249;
			{8'd33, 8'd118}: color_data = 12'h249;
			{8'd33, 8'd119}: color_data = 12'h249;
			{8'd33, 8'd120}: color_data = 12'h249;
			{8'd33, 8'd121}: color_data = 12'h249;
			{8'd33, 8'd122}: color_data = 12'h136;
			{8'd33, 8'd123}: color_data = 12'h000;
			{8'd33, 8'd136}: color_data = 12'h000;
			{8'd33, 8'd137}: color_data = 12'h321;
			{8'd33, 8'd138}: color_data = 12'h532;
			{8'd33, 8'd139}: color_data = 12'h633;
			{8'd33, 8'd140}: color_data = 12'h432;
			{8'd33, 8'd141}: color_data = 12'h111;
			{8'd33, 8'd142}: color_data = 12'h000;
			{8'd34, 8'd17}: color_data = 12'hfc5;
			{8'd34, 8'd18}: color_data = 12'hfc5;
			{8'd34, 8'd19}: color_data = 12'hfc4;
			{8'd34, 8'd20}: color_data = 12'hd90;
			{8'd34, 8'd21}: color_data = 12'hd90;
			{8'd34, 8'd22}: color_data = 12'hd90;
			{8'd34, 8'd23}: color_data = 12'hd90;
			{8'd34, 8'd24}: color_data = 12'hea1;
			{8'd34, 8'd25}: color_data = 12'heb2;
			{8'd34, 8'd26}: color_data = 12'hd90;
			{8'd34, 8'd27}: color_data = 12'hd90;
			{8'd34, 8'd28}: color_data = 12'hd90;
			{8'd34, 8'd29}: color_data = 12'hd90;
			{8'd34, 8'd30}: color_data = 12'hea0;
			{8'd34, 8'd31}: color_data = 12'hfc4;
			{8'd34, 8'd32}: color_data = 12'heb3;
			{8'd34, 8'd33}: color_data = 12'heb2;
			{8'd34, 8'd34}: color_data = 12'hfc5;
			{8'd34, 8'd35}: color_data = 12'hfc4;
			{8'd34, 8'd36}: color_data = 12'hfa5;
			{8'd34, 8'd54}: color_data = 12'h000;
			{8'd34, 8'd55}: color_data = 12'h000;
			{8'd34, 8'd56}: color_data = 12'h000;
			{8'd34, 8'd57}: color_data = 12'h000;
			{8'd34, 8'd58}: color_data = 12'h000;
			{8'd34, 8'd59}: color_data = 12'h000;
			{8'd34, 8'd60}: color_data = 12'h000;
			{8'd34, 8'd61}: color_data = 12'h000;
			{8'd34, 8'd62}: color_data = 12'h051;
			{8'd34, 8'd63}: color_data = 12'h0a3;
			{8'd34, 8'd64}: color_data = 12'h0a3;
			{8'd34, 8'd65}: color_data = 12'h0a3;
			{8'd34, 8'd66}: color_data = 12'h0a3;
			{8'd34, 8'd67}: color_data = 12'h0a3;
			{8'd34, 8'd68}: color_data = 12'h062;
			{8'd34, 8'd69}: color_data = 12'hca9;
			{8'd34, 8'd70}: color_data = 12'hfdb;
			{8'd34, 8'd71}: color_data = 12'heca;
			{8'd34, 8'd72}: color_data = 12'h876;
			{8'd34, 8'd73}: color_data = 12'hb98;
			{8'd34, 8'd74}: color_data = 12'hfda;
			{8'd34, 8'd75}: color_data = 12'h332;
			{8'd34, 8'd76}: color_data = 12'hba8;
			{8'd34, 8'd77}: color_data = 12'hb98;
			{8'd34, 8'd78}: color_data = 12'hfdb;
			{8'd34, 8'd79}: color_data = 12'hfdb;
			{8'd34, 8'd80}: color_data = 12'hfeb;
			{8'd34, 8'd81}: color_data = 12'h765;
			{8'd34, 8'd82}: color_data = 12'h000;
			{8'd34, 8'd83}: color_data = 12'h000;
			{8'd34, 8'd84}: color_data = 12'h543;
			{8'd34, 8'd85}: color_data = 12'hfdb;
			{8'd34, 8'd86}: color_data = 12'hfdb;
			{8'd34, 8'd87}: color_data = 12'hfdb;
			{8'd34, 8'd88}: color_data = 12'hfdb;
			{8'd34, 8'd89}: color_data = 12'ha97;
			{8'd34, 8'd90}: color_data = 12'heca;
			{8'd34, 8'd91}: color_data = 12'hfeb;
			{8'd34, 8'd92}: color_data = 12'ha98;
			{8'd34, 8'd93}: color_data = 12'h083;
			{8'd34, 8'd94}: color_data = 12'h0a3;
			{8'd34, 8'd95}: color_data = 12'h0a3;
			{8'd34, 8'd96}: color_data = 12'h0a3;
			{8'd34, 8'd97}: color_data = 12'h0a3;
			{8'd34, 8'd98}: color_data = 12'h082;
			{8'd34, 8'd99}: color_data = 12'h586;
			{8'd34, 8'd100}: color_data = 12'h274;
			{8'd34, 8'd101}: color_data = 12'h083;
			{8'd34, 8'd102}: color_data = 12'h052;
			{8'd34, 8'd103}: color_data = 12'h024;
			{8'd34, 8'd104}: color_data = 12'h136;
			{8'd34, 8'd105}: color_data = 12'h136;
			{8'd34, 8'd106}: color_data = 12'h136;
			{8'd34, 8'd107}: color_data = 12'h136;
			{8'd34, 8'd108}: color_data = 12'h137;
			{8'd34, 8'd109}: color_data = 12'h249;
			{8'd34, 8'd110}: color_data = 12'h249;
			{8'd34, 8'd111}: color_data = 12'h249;
			{8'd34, 8'd112}: color_data = 12'h249;
			{8'd34, 8'd113}: color_data = 12'h249;
			{8'd34, 8'd114}: color_data = 12'h249;
			{8'd34, 8'd115}: color_data = 12'h249;
			{8'd34, 8'd116}: color_data = 12'h249;
			{8'd34, 8'd117}: color_data = 12'h249;
			{8'd34, 8'd118}: color_data = 12'h249;
			{8'd34, 8'd119}: color_data = 12'h249;
			{8'd34, 8'd120}: color_data = 12'h249;
			{8'd34, 8'd121}: color_data = 12'h249;
			{8'd34, 8'd122}: color_data = 12'h013;
			{8'd34, 8'd137}: color_data = 12'h000;
			{8'd34, 8'd138}: color_data = 12'h100;
			{8'd34, 8'd139}: color_data = 12'h110;
			{8'd34, 8'd140}: color_data = 12'h000;
			{8'd34, 8'd141}: color_data = 12'h000;
			{8'd35, 8'd17}: color_data = 12'hfc5;
			{8'd35, 8'd18}: color_data = 12'hfc5;
			{8'd35, 8'd19}: color_data = 12'hfc5;
			{8'd35, 8'd20}: color_data = 12'hea1;
			{8'd35, 8'd21}: color_data = 12'hd90;
			{8'd35, 8'd22}: color_data = 12'hd90;
			{8'd35, 8'd23}: color_data = 12'hd90;
			{8'd35, 8'd24}: color_data = 12'hd90;
			{8'd35, 8'd25}: color_data = 12'hd90;
			{8'd35, 8'd26}: color_data = 12'hd90;
			{8'd35, 8'd27}: color_data = 12'hd90;
			{8'd35, 8'd28}: color_data = 12'hd90;
			{8'd35, 8'd29}: color_data = 12'hd90;
			{8'd35, 8'd30}: color_data = 12'hd90;
			{8'd35, 8'd31}: color_data = 12'hfb3;
			{8'd35, 8'd32}: color_data = 12'hfc6;
			{8'd35, 8'd33}: color_data = 12'hfc5;
			{8'd35, 8'd34}: color_data = 12'hfc5;
			{8'd35, 8'd35}: color_data = 12'hfc5;
			{8'd35, 8'd61}: color_data = 12'h041;
			{8'd35, 8'd62}: color_data = 12'h0a3;
			{8'd35, 8'd63}: color_data = 12'h0a3;
			{8'd35, 8'd64}: color_data = 12'h0a3;
			{8'd35, 8'd65}: color_data = 12'h0a3;
			{8'd35, 8'd66}: color_data = 12'h0a3;
			{8'd35, 8'd67}: color_data = 12'h062;
			{8'd35, 8'd68}: color_data = 12'h321;
			{8'd35, 8'd69}: color_data = 12'hdb9;
			{8'd35, 8'd70}: color_data = 12'hfeb;
			{8'd35, 8'd71}: color_data = 12'hfdb;
			{8'd35, 8'd72}: color_data = 12'hfdb;
			{8'd35, 8'd73}: color_data = 12'h554;
			{8'd35, 8'd74}: color_data = 12'ha97;
			{8'd35, 8'd75}: color_data = 12'h433;
			{8'd35, 8'd76}: color_data = 12'ha87;
			{8'd35, 8'd77}: color_data = 12'hfda;
			{8'd35, 8'd78}: color_data = 12'hfdb;
			{8'd35, 8'd79}: color_data = 12'hfdb;
			{8'd35, 8'd80}: color_data = 12'hfdb;
			{8'd35, 8'd81}: color_data = 12'ha97;
			{8'd35, 8'd82}: color_data = 12'h000;
			{8'd35, 8'd83}: color_data = 12'h000;
			{8'd35, 8'd84}: color_data = 12'h322;
			{8'd35, 8'd85}: color_data = 12'hfdb;
			{8'd35, 8'd86}: color_data = 12'hfdb;
			{8'd35, 8'd87}: color_data = 12'hfdb;
			{8'd35, 8'd88}: color_data = 12'hfdb;
			{8'd35, 8'd89}: color_data = 12'ha97;
			{8'd35, 8'd90}: color_data = 12'hfdb;
			{8'd35, 8'd91}: color_data = 12'hfdb;
			{8'd35, 8'd92}: color_data = 12'h574;
			{8'd35, 8'd93}: color_data = 12'h0a3;
			{8'd35, 8'd94}: color_data = 12'h0a3;
			{8'd35, 8'd95}: color_data = 12'h083;
			{8'd35, 8'd96}: color_data = 12'h274;
			{8'd35, 8'd97}: color_data = 12'h586;
			{8'd35, 8'd98}: color_data = 12'haaa;
			{8'd35, 8'd99}: color_data = 12'hfff;
			{8'd35, 8'd100}: color_data = 12'hddd;
			{8'd35, 8'd101}: color_data = 12'hddd;
			{8'd35, 8'd102}: color_data = 12'hddd;
			{8'd35, 8'd103}: color_data = 12'h778;
			{8'd35, 8'd104}: color_data = 12'h346;
			{8'd35, 8'd105}: color_data = 12'h236;
			{8'd35, 8'd106}: color_data = 12'h236;
			{8'd35, 8'd107}: color_data = 12'h137;
			{8'd35, 8'd108}: color_data = 12'h137;
			{8'd35, 8'd109}: color_data = 12'h125;
			{8'd35, 8'd110}: color_data = 12'h248;
			{8'd35, 8'd111}: color_data = 12'h249;
			{8'd35, 8'd112}: color_data = 12'h249;
			{8'd35, 8'd113}: color_data = 12'h249;
			{8'd35, 8'd114}: color_data = 12'h249;
			{8'd35, 8'd115}: color_data = 12'h249;
			{8'd35, 8'd116}: color_data = 12'h249;
			{8'd35, 8'd117}: color_data = 12'h249;
			{8'd35, 8'd118}: color_data = 12'h249;
			{8'd35, 8'd119}: color_data = 12'h249;
			{8'd35, 8'd120}: color_data = 12'h249;
			{8'd35, 8'd121}: color_data = 12'h136;
			{8'd35, 8'd122}: color_data = 12'h000;
			{8'd36, 8'd18}: color_data = 12'hfc5;
			{8'd36, 8'd19}: color_data = 12'hfc5;
			{8'd36, 8'd20}: color_data = 12'heb2;
			{8'd36, 8'd21}: color_data = 12'hd90;
			{8'd36, 8'd22}: color_data = 12'hd90;
			{8'd36, 8'd23}: color_data = 12'hd90;
			{8'd36, 8'd24}: color_data = 12'hd90;
			{8'd36, 8'd25}: color_data = 12'hd90;
			{8'd36, 8'd26}: color_data = 12'hd90;
			{8'd36, 8'd27}: color_data = 12'hd90;
			{8'd36, 8'd28}: color_data = 12'hd90;
			{8'd36, 8'd29}: color_data = 12'hd90;
			{8'd36, 8'd30}: color_data = 12'hd90;
			{8'd36, 8'd31}: color_data = 12'hea1;
			{8'd36, 8'd32}: color_data = 12'hfc5;
			{8'd36, 8'd33}: color_data = 12'hfc5;
			{8'd36, 8'd34}: color_data = 12'hfc5;
			{8'd36, 8'd35}: color_data = 12'hfc5;
			{8'd36, 8'd60}: color_data = 12'h010;
			{8'd36, 8'd61}: color_data = 12'h083;
			{8'd36, 8'd62}: color_data = 12'h0a3;
			{8'd36, 8'd63}: color_data = 12'h0a3;
			{8'd36, 8'd64}: color_data = 12'h0a3;
			{8'd36, 8'd65}: color_data = 12'h0a3;
			{8'd36, 8'd66}: color_data = 12'h062;
			{8'd36, 8'd67}: color_data = 12'h421;
			{8'd36, 8'd68}: color_data = 12'h742;
			{8'd36, 8'd69}: color_data = 12'h532;
			{8'd36, 8'd70}: color_data = 12'hdb9;
			{8'd36, 8'd71}: color_data = 12'hfec;
			{8'd36, 8'd72}: color_data = 12'h654;
			{8'd36, 8'd73}: color_data = 12'h765;
			{8'd36, 8'd74}: color_data = 12'ha87;
			{8'd36, 8'd75}: color_data = 12'hca9;
			{8'd36, 8'd76}: color_data = 12'hfeb;
			{8'd36, 8'd77}: color_data = 12'hfdb;
			{8'd36, 8'd78}: color_data = 12'hfdb;
			{8'd36, 8'd79}: color_data = 12'hfdb;
			{8'd36, 8'd80}: color_data = 12'hfdb;
			{8'd36, 8'd81}: color_data = 12'hfeb;
			{8'd36, 8'd82}: color_data = 12'h543;
			{8'd36, 8'd83}: color_data = 12'h000;
			{8'd36, 8'd84}: color_data = 12'h876;
			{8'd36, 8'd85}: color_data = 12'hfeb;
			{8'd36, 8'd86}: color_data = 12'hfdb;
			{8'd36, 8'd87}: color_data = 12'hfdb;
			{8'd36, 8'd88}: color_data = 12'hfdb;
			{8'd36, 8'd89}: color_data = 12'h986;
			{8'd36, 8'd90}: color_data = 12'hba8;
			{8'd36, 8'd91}: color_data = 12'h886;
			{8'd36, 8'd92}: color_data = 12'h083;
			{8'd36, 8'd93}: color_data = 12'h0b3;
			{8'd36, 8'd94}: color_data = 12'h173;
			{8'd36, 8'd95}: color_data = 12'hbbb;
			{8'd36, 8'd96}: color_data = 12'hfff;
			{8'd36, 8'd97}: color_data = 12'hfff;
			{8'd36, 8'd98}: color_data = 12'hfff;
			{8'd36, 8'd99}: color_data = 12'hfff;
			{8'd36, 8'd100}: color_data = 12'hfff;
			{8'd36, 8'd101}: color_data = 12'hfff;
			{8'd36, 8'd102}: color_data = 12'hfff;
			{8'd36, 8'd103}: color_data = 12'hfff;
			{8'd36, 8'd104}: color_data = 12'hfff;
			{8'd36, 8'd105}: color_data = 12'haa8;
			{8'd36, 8'd106}: color_data = 12'hcb0;
			{8'd36, 8'd107}: color_data = 12'haa0;
			{8'd36, 8'd108}: color_data = 12'h247;
			{8'd36, 8'd109}: color_data = 12'h248;
			{8'd36, 8'd110}: color_data = 12'h135;
			{8'd36, 8'd111}: color_data = 12'h249;
			{8'd36, 8'd112}: color_data = 12'h249;
			{8'd36, 8'd113}: color_data = 12'h249;
			{8'd36, 8'd114}: color_data = 12'h249;
			{8'd36, 8'd115}: color_data = 12'h249;
			{8'd36, 8'd116}: color_data = 12'h249;
			{8'd36, 8'd117}: color_data = 12'h249;
			{8'd36, 8'd118}: color_data = 12'h249;
			{8'd36, 8'd119}: color_data = 12'h249;
			{8'd36, 8'd120}: color_data = 12'h249;
			{8'd36, 8'd121}: color_data = 12'h124;
			{8'd37, 8'd18}: color_data = 12'hfc6;
			{8'd37, 8'd19}: color_data = 12'hfc5;
			{8'd37, 8'd20}: color_data = 12'hfc4;
			{8'd37, 8'd21}: color_data = 12'hda0;
			{8'd37, 8'd22}: color_data = 12'hd90;
			{8'd37, 8'd23}: color_data = 12'hd90;
			{8'd37, 8'd24}: color_data = 12'hd90;
			{8'd37, 8'd25}: color_data = 12'hd90;
			{8'd37, 8'd26}: color_data = 12'hd90;
			{8'd37, 8'd27}: color_data = 12'hd90;
			{8'd37, 8'd28}: color_data = 12'hd90;
			{8'd37, 8'd29}: color_data = 12'hd90;
			{8'd37, 8'd30}: color_data = 12'hd90;
			{8'd37, 8'd31}: color_data = 12'hd90;
			{8'd37, 8'd32}: color_data = 12'heb3;
			{8'd37, 8'd33}: color_data = 12'hfc5;
			{8'd37, 8'd34}: color_data = 12'hfc6;
			{8'd37, 8'd59}: color_data = 12'h000;
			{8'd37, 8'd60}: color_data = 12'h051;
			{8'd37, 8'd61}: color_data = 12'h0a3;
			{8'd37, 8'd62}: color_data = 12'h0a3;
			{8'd37, 8'd63}: color_data = 12'h0a3;
			{8'd37, 8'd64}: color_data = 12'h0a3;
			{8'd37, 8'd65}: color_data = 12'h052;
			{8'd37, 8'd66}: color_data = 12'h000;
			{8'd37, 8'd67}: color_data = 12'h000;
			{8'd37, 8'd68}: color_data = 12'h210;
			{8'd37, 8'd69}: color_data = 12'h100;
			{8'd37, 8'd70}: color_data = 12'h211;
			{8'd37, 8'd71}: color_data = 12'h986;
			{8'd37, 8'd72}: color_data = 12'h554;
			{8'd37, 8'd73}: color_data = 12'h765;
			{8'd37, 8'd74}: color_data = 12'hb98;
			{8'd37, 8'd75}: color_data = 12'hfeb;
			{8'd37, 8'd76}: color_data = 12'hfdb;
			{8'd37, 8'd77}: color_data = 12'hfdb;
			{8'd37, 8'd78}: color_data = 12'hfdb;
			{8'd37, 8'd79}: color_data = 12'hfdb;
			{8'd37, 8'd80}: color_data = 12'hfdb;
			{8'd37, 8'd81}: color_data = 12'hfeb;
			{8'd37, 8'd82}: color_data = 12'ha97;
			{8'd37, 8'd83}: color_data = 12'h000;
			{8'd37, 8'd84}: color_data = 12'hca9;
			{8'd37, 8'd85}: color_data = 12'hfeb;
			{8'd37, 8'd86}: color_data = 12'hfdb;
			{8'd37, 8'd87}: color_data = 12'hfdb;
			{8'd37, 8'd88}: color_data = 12'hfdb;
			{8'd37, 8'd89}: color_data = 12'h566;
			{8'd37, 8'd90}: color_data = 12'h043;
			{8'd37, 8'd91}: color_data = 12'h082;
			{8'd37, 8'd92}: color_data = 12'h093;
			{8'd37, 8'd93}: color_data = 12'h062;
			{8'd37, 8'd94}: color_data = 12'h566;
			{8'd37, 8'd95}: color_data = 12'hfff;
			{8'd37, 8'd96}: color_data = 12'hfff;
			{8'd37, 8'd97}: color_data = 12'hfff;
			{8'd37, 8'd98}: color_data = 12'hfff;
			{8'd37, 8'd99}: color_data = 12'hfff;
			{8'd37, 8'd100}: color_data = 12'hfff;
			{8'd37, 8'd101}: color_data = 12'hfff;
			{8'd37, 8'd102}: color_data = 12'hfff;
			{8'd37, 8'd103}: color_data = 12'hfff;
			{8'd37, 8'd104}: color_data = 12'hfff;
			{8'd37, 8'd105}: color_data = 12'hddd;
			{8'd37, 8'd106}: color_data = 12'hcc0;
			{8'd37, 8'd107}: color_data = 12'hdd0;
			{8'd37, 8'd108}: color_data = 12'h236;
			{8'd37, 8'd109}: color_data = 12'h137;
			{8'd37, 8'd110}: color_data = 12'h136;
			{8'd37, 8'd111}: color_data = 12'h249;
			{8'd37, 8'd112}: color_data = 12'h249;
			{8'd37, 8'd113}: color_data = 12'h249;
			{8'd37, 8'd114}: color_data = 12'h249;
			{8'd37, 8'd115}: color_data = 12'h249;
			{8'd37, 8'd116}: color_data = 12'h249;
			{8'd37, 8'd117}: color_data = 12'h249;
			{8'd37, 8'd118}: color_data = 12'h249;
			{8'd37, 8'd119}: color_data = 12'h249;
			{8'd37, 8'd120}: color_data = 12'h248;
			{8'd37, 8'd121}: color_data = 12'h001;
			{8'd38, 8'd17}: color_data = 12'hfc4;
			{8'd38, 8'd18}: color_data = 12'hfc5;
			{8'd38, 8'd19}: color_data = 12'hfc5;
			{8'd38, 8'd20}: color_data = 12'hfc5;
			{8'd38, 8'd21}: color_data = 12'hfc4;
			{8'd38, 8'd22}: color_data = 12'hea1;
			{8'd38, 8'd23}: color_data = 12'hda0;
			{8'd38, 8'd24}: color_data = 12'hd90;
			{8'd38, 8'd25}: color_data = 12'hd90;
			{8'd38, 8'd26}: color_data = 12'hd90;
			{8'd38, 8'd27}: color_data = 12'heb2;
			{8'd38, 8'd28}: color_data = 12'heb2;
			{8'd38, 8'd29}: color_data = 12'hd90;
			{8'd38, 8'd30}: color_data = 12'hd90;
			{8'd38, 8'd31}: color_data = 12'hd90;
			{8'd38, 8'd32}: color_data = 12'hea1;
			{8'd38, 8'd33}: color_data = 12'hfc5;
			{8'd38, 8'd34}: color_data = 12'hfc5;
			{8'd38, 8'd35}: color_data = 12'hfc5;
			{8'd38, 8'd59}: color_data = 12'h000;
			{8'd38, 8'd60}: color_data = 12'h082;
			{8'd38, 8'd61}: color_data = 12'h0a4;
			{8'd38, 8'd62}: color_data = 12'h0a4;
			{8'd38, 8'd63}: color_data = 12'h093;
			{8'd38, 8'd64}: color_data = 12'h041;
			{8'd38, 8'd65}: color_data = 12'h000;
			{8'd38, 8'd71}: color_data = 12'h221;
			{8'd38, 8'd72}: color_data = 12'h876;
			{8'd38, 8'd73}: color_data = 12'h543;
			{8'd38, 8'd74}: color_data = 12'hfdb;
			{8'd38, 8'd75}: color_data = 12'hfdb;
			{8'd38, 8'd76}: color_data = 12'hfdb;
			{8'd38, 8'd77}: color_data = 12'hfdb;
			{8'd38, 8'd78}: color_data = 12'hfdb;
			{8'd38, 8'd79}: color_data = 12'hfdb;
			{8'd38, 8'd80}: color_data = 12'hfdb;
			{8'd38, 8'd81}: color_data = 12'hfeb;
			{8'd38, 8'd82}: color_data = 12'hb98;
			{8'd38, 8'd83}: color_data = 12'h000;
			{8'd38, 8'd84}: color_data = 12'ha87;
			{8'd38, 8'd85}: color_data = 12'heca;
			{8'd38, 8'd86}: color_data = 12'hfdb;
			{8'd38, 8'd87}: color_data = 12'hfeb;
			{8'd38, 8'd88}: color_data = 12'hdb9;
			{8'd38, 8'd89}: color_data = 12'h468;
			{8'd38, 8'd90}: color_data = 12'h479;
			{8'd38, 8'd91}: color_data = 12'h043;
			{8'd38, 8'd92}: color_data = 12'h136;
			{8'd38, 8'd93}: color_data = 12'h137;
			{8'd38, 8'd94}: color_data = 12'h446;
			{8'd38, 8'd95}: color_data = 12'hfff;
			{8'd38, 8'd96}: color_data = 12'hfff;
			{8'd38, 8'd97}: color_data = 12'hfff;
			{8'd38, 8'd98}: color_data = 12'hfff;
			{8'd38, 8'd99}: color_data = 12'hfff;
			{8'd38, 8'd100}: color_data = 12'hfff;
			{8'd38, 8'd101}: color_data = 12'hfff;
			{8'd38, 8'd102}: color_data = 12'hfff;
			{8'd38, 8'd103}: color_data = 12'hfff;
			{8'd38, 8'd104}: color_data = 12'hfff;
			{8'd38, 8'd105}: color_data = 12'heee;
			{8'd38, 8'd106}: color_data = 12'h552;
			{8'd38, 8'd107}: color_data = 12'h232;
			{8'd38, 8'd108}: color_data = 12'h125;
			{8'd38, 8'd109}: color_data = 12'h136;
			{8'd38, 8'd110}: color_data = 12'h249;
			{8'd38, 8'd111}: color_data = 12'h249;
			{8'd38, 8'd112}: color_data = 12'h249;
			{8'd38, 8'd113}: color_data = 12'h249;
			{8'd38, 8'd114}: color_data = 12'h249;
			{8'd38, 8'd115}: color_data = 12'h249;
			{8'd38, 8'd116}: color_data = 12'h249;
			{8'd38, 8'd117}: color_data = 12'h249;
			{8'd38, 8'd118}: color_data = 12'h249;
			{8'd38, 8'd119}: color_data = 12'h249;
			{8'd38, 8'd120}: color_data = 12'h136;
			{8'd38, 8'd121}: color_data = 12'h000;
			{8'd39, 8'd16}: color_data = 12'hfc5;
			{8'd39, 8'd17}: color_data = 12'hfc4;
			{8'd39, 8'd18}: color_data = 12'hfc5;
			{8'd39, 8'd19}: color_data = 12'hfc5;
			{8'd39, 8'd20}: color_data = 12'hfc5;
			{8'd39, 8'd21}: color_data = 12'hfc6;
			{8'd39, 8'd22}: color_data = 12'hfc6;
			{8'd39, 8'd23}: color_data = 12'hfc5;
			{8'd39, 8'd24}: color_data = 12'hfc4;
			{8'd39, 8'd25}: color_data = 12'hfb3;
			{8'd39, 8'd26}: color_data = 12'hfc4;
			{8'd39, 8'd27}: color_data = 12'hfc5;
			{8'd39, 8'd28}: color_data = 12'hfc5;
			{8'd39, 8'd29}: color_data = 12'hda0;
			{8'd39, 8'd30}: color_data = 12'hd90;
			{8'd39, 8'd31}: color_data = 12'hd90;
			{8'd39, 8'd32}: color_data = 12'hfb3;
			{8'd39, 8'd33}: color_data = 12'hfc5;
			{8'd39, 8'd34}: color_data = 12'hfc5;
			{8'd39, 8'd35}: color_data = 12'hfb7;
			{8'd39, 8'd59}: color_data = 12'h000;
			{8'd39, 8'd60}: color_data = 12'h062;
			{8'd39, 8'd61}: color_data = 12'h093;
			{8'd39, 8'd62}: color_data = 12'h062;
			{8'd39, 8'd63}: color_data = 12'h021;
			{8'd39, 8'd64}: color_data = 12'h000;
			{8'd39, 8'd71}: color_data = 12'h210;
			{8'd39, 8'd72}: color_data = 12'h653;
			{8'd39, 8'd73}: color_data = 12'h986;
			{8'd39, 8'd74}: color_data = 12'hfdb;
			{8'd39, 8'd75}: color_data = 12'hfdb;
			{8'd39, 8'd76}: color_data = 12'hfdb;
			{8'd39, 8'd77}: color_data = 12'hfdb;
			{8'd39, 8'd78}: color_data = 12'hfdb;
			{8'd39, 8'd79}: color_data = 12'hfdb;
			{8'd39, 8'd80}: color_data = 12'hfdb;
			{8'd39, 8'd81}: color_data = 12'hfeb;
			{8'd39, 8'd82}: color_data = 12'h876;
			{8'd39, 8'd83}: color_data = 12'h000;
			{8'd39, 8'd84}: color_data = 12'ha87;
			{8'd39, 8'd85}: color_data = 12'hca8;
			{8'd39, 8'd86}: color_data = 12'hfec;
			{8'd39, 8'd87}: color_data = 12'heca;
			{8'd39, 8'd88}: color_data = 12'h566;
			{8'd39, 8'd89}: color_data = 12'h48a;
			{8'd39, 8'd90}: color_data = 12'h59b;
			{8'd39, 8'd91}: color_data = 12'h368;
			{8'd39, 8'd92}: color_data = 12'h125;
			{8'd39, 8'd93}: color_data = 12'h257;
			{8'd39, 8'd94}: color_data = 12'h367;
			{8'd39, 8'd95}: color_data = 12'hddd;
			{8'd39, 8'd96}: color_data = 12'hfff;
			{8'd39, 8'd97}: color_data = 12'hfff;
			{8'd39, 8'd98}: color_data = 12'hfff;
			{8'd39, 8'd99}: color_data = 12'hfff;
			{8'd39, 8'd100}: color_data = 12'hfff;
			{8'd39, 8'd101}: color_data = 12'hfff;
			{8'd39, 8'd102}: color_data = 12'heee;
			{8'd39, 8'd103}: color_data = 12'hfff;
			{8'd39, 8'd104}: color_data = 12'hfff;
			{8'd39, 8'd105}: color_data = 12'hffe;
			{8'd39, 8'd106}: color_data = 12'h235;
			{8'd39, 8'd107}: color_data = 12'h137;
			{8'd39, 8'd108}: color_data = 12'h249;
			{8'd39, 8'd109}: color_data = 12'h249;
			{8'd39, 8'd110}: color_data = 12'h249;
			{8'd39, 8'd111}: color_data = 12'h249;
			{8'd39, 8'd112}: color_data = 12'h249;
			{8'd39, 8'd113}: color_data = 12'h249;
			{8'd39, 8'd114}: color_data = 12'h249;
			{8'd39, 8'd115}: color_data = 12'h249;
			{8'd39, 8'd116}: color_data = 12'h249;
			{8'd39, 8'd117}: color_data = 12'h249;
			{8'd39, 8'd118}: color_data = 12'h249;
			{8'd39, 8'd119}: color_data = 12'h249;
			{8'd39, 8'd120}: color_data = 12'h136;
			{8'd39, 8'd121}: color_data = 12'h000;
			{8'd40, 8'd16}: color_data = 12'hfc4;
			{8'd40, 8'd17}: color_data = 12'hfc5;
			{8'd40, 8'd18}: color_data = 12'hfb3;
			{8'd40, 8'd19}: color_data = 12'hea1;
			{8'd40, 8'd20}: color_data = 12'hea2;
			{8'd40, 8'd21}: color_data = 12'hea1;
			{8'd40, 8'd22}: color_data = 12'hea1;
			{8'd40, 8'd23}: color_data = 12'heb2;
			{8'd40, 8'd24}: color_data = 12'hfb4;
			{8'd40, 8'd25}: color_data = 12'hfc5;
			{8'd40, 8'd26}: color_data = 12'hfc6;
			{8'd40, 8'd27}: color_data = 12'hfc5;
			{8'd40, 8'd28}: color_data = 12'hfc6;
			{8'd40, 8'd29}: color_data = 12'heb3;
			{8'd40, 8'd30}: color_data = 12'hd90;
			{8'd40, 8'd31}: color_data = 12'heb2;
			{8'd40, 8'd32}: color_data = 12'hfc5;
			{8'd40, 8'd33}: color_data = 12'hfc4;
			{8'd40, 8'd34}: color_data = 12'hec5;
			{8'd40, 8'd60}: color_data = 12'h010;
			{8'd40, 8'd61}: color_data = 12'h010;
			{8'd40, 8'd62}: color_data = 12'h000;
			{8'd40, 8'd70}: color_data = 12'h000;
			{8'd40, 8'd71}: color_data = 12'h873;
			{8'd40, 8'd72}: color_data = 12'hca5;
			{8'd40, 8'd73}: color_data = 12'hb97;
			{8'd40, 8'd74}: color_data = 12'hfdb;
			{8'd40, 8'd75}: color_data = 12'hfdb;
			{8'd40, 8'd76}: color_data = 12'hfdb;
			{8'd40, 8'd77}: color_data = 12'hfdb;
			{8'd40, 8'd78}: color_data = 12'hfdb;
			{8'd40, 8'd79}: color_data = 12'hfdb;
			{8'd40, 8'd80}: color_data = 12'hfdb;
			{8'd40, 8'd81}: color_data = 12'hfdb;
			{8'd40, 8'd82}: color_data = 12'h765;
			{8'd40, 8'd83}: color_data = 12'hba8;
			{8'd40, 8'd84}: color_data = 12'ha87;
			{8'd40, 8'd85}: color_data = 12'ha97;
			{8'd40, 8'd86}: color_data = 12'h766;
			{8'd40, 8'd87}: color_data = 12'h122;
			{8'd40, 8'd88}: color_data = 12'h379;
			{8'd40, 8'd89}: color_data = 12'h49b;
			{8'd40, 8'd90}: color_data = 12'h48a;
			{8'd40, 8'd91}: color_data = 12'h256;
			{8'd40, 8'd92}: color_data = 12'h378;
			{8'd40, 8'd93}: color_data = 12'h59b;
			{8'd40, 8'd94}: color_data = 12'h368;
			{8'd40, 8'd95}: color_data = 12'haaa;
			{8'd40, 8'd96}: color_data = 12'hfff;
			{8'd40, 8'd97}: color_data = 12'hfff;
			{8'd40, 8'd98}: color_data = 12'hfff;
			{8'd40, 8'd99}: color_data = 12'heee;
			{8'd40, 8'd100}: color_data = 12'hbbb;
			{8'd40, 8'd101}: color_data = 12'hfff;
			{8'd40, 8'd102}: color_data = 12'haaa;
			{8'd40, 8'd103}: color_data = 12'hfff;
			{8'd40, 8'd104}: color_data = 12'hfff;
			{8'd40, 8'd105}: color_data = 12'heee;
			{8'd40, 8'd106}: color_data = 12'h556;
			{8'd40, 8'd107}: color_data = 12'h247;
			{8'd40, 8'd108}: color_data = 12'h249;
			{8'd40, 8'd109}: color_data = 12'h249;
			{8'd40, 8'd110}: color_data = 12'h249;
			{8'd40, 8'd111}: color_data = 12'h249;
			{8'd40, 8'd112}: color_data = 12'h249;
			{8'd40, 8'd113}: color_data = 12'h249;
			{8'd40, 8'd114}: color_data = 12'h249;
			{8'd40, 8'd115}: color_data = 12'h249;
			{8'd40, 8'd116}: color_data = 12'h249;
			{8'd40, 8'd117}: color_data = 12'h249;
			{8'd40, 8'd118}: color_data = 12'h249;
			{8'd40, 8'd119}: color_data = 12'h249;
			{8'd40, 8'd120}: color_data = 12'h137;
			{8'd40, 8'd121}: color_data = 12'h000;
			{8'd40, 8'd129}: color_data = 12'h000;
			{8'd40, 8'd130}: color_data = 12'h000;
			{8'd40, 8'd131}: color_data = 12'h000;
			{8'd40, 8'd132}: color_data = 12'h211;
			{8'd40, 8'd133}: color_data = 12'h311;
			{8'd40, 8'd134}: color_data = 12'h211;
			{8'd40, 8'd135}: color_data = 12'h000;
			{8'd41, 8'd15}: color_data = 12'hfc3;
			{8'd41, 8'd16}: color_data = 12'hfc4;
			{8'd41, 8'd17}: color_data = 12'hfc5;
			{8'd41, 8'd18}: color_data = 12'hda0;
			{8'd41, 8'd19}: color_data = 12'hd90;
			{8'd41, 8'd20}: color_data = 12'hd90;
			{8'd41, 8'd21}: color_data = 12'hd90;
			{8'd41, 8'd22}: color_data = 12'hd90;
			{8'd41, 8'd23}: color_data = 12'hd90;
			{8'd41, 8'd24}: color_data = 12'hd90;
			{8'd41, 8'd25}: color_data = 12'hda0;
			{8'd41, 8'd26}: color_data = 12'hea2;
			{8'd41, 8'd27}: color_data = 12'hfb3;
			{8'd41, 8'd28}: color_data = 12'hfc5;
			{8'd41, 8'd29}: color_data = 12'hfc5;
			{8'd41, 8'd30}: color_data = 12'heb2;
			{8'd41, 8'd31}: color_data = 12'hfc5;
			{8'd41, 8'd32}: color_data = 12'hfc5;
			{8'd41, 8'd33}: color_data = 12'hfc5;
			{8'd41, 8'd68}: color_data = 12'h000;
			{8'd41, 8'd69}: color_data = 12'h221;
			{8'd41, 8'd70}: color_data = 12'h663;
			{8'd41, 8'd71}: color_data = 12'h873;
			{8'd41, 8'd72}: color_data = 12'ha84;
			{8'd41, 8'd73}: color_data = 12'ha97;
			{8'd41, 8'd74}: color_data = 12'hfeb;
			{8'd41, 8'd75}: color_data = 12'hfdb;
			{8'd41, 8'd76}: color_data = 12'hfdb;
			{8'd41, 8'd77}: color_data = 12'hfdb;
			{8'd41, 8'd78}: color_data = 12'hfdb;
			{8'd41, 8'd79}: color_data = 12'hfdb;
			{8'd41, 8'd80}: color_data = 12'hfeb;
			{8'd41, 8'd81}: color_data = 12'hb98;
			{8'd41, 8'd82}: color_data = 12'hcb9;
			{8'd41, 8'd83}: color_data = 12'hfda;
			{8'd41, 8'd84}: color_data = 12'h456;
			{8'd41, 8'd85}: color_data = 12'h256;
			{8'd41, 8'd86}: color_data = 12'h001;
			{8'd41, 8'd87}: color_data = 12'h123;
			{8'd41, 8'd88}: color_data = 12'h48a;
			{8'd41, 8'd89}: color_data = 12'h49b;
			{8'd41, 8'd90}: color_data = 12'h367;
			{8'd41, 8'd91}: color_data = 12'h378;
			{8'd41, 8'd92}: color_data = 12'h59b;
			{8'd41, 8'd93}: color_data = 12'h367;
			{8'd41, 8'd94}: color_data = 12'h062;
			{8'd41, 8'd95}: color_data = 12'h586;
			{8'd41, 8'd96}: color_data = 12'hfff;
			{8'd41, 8'd97}: color_data = 12'heee;
			{8'd41, 8'd98}: color_data = 12'haaa;
			{8'd41, 8'd99}: color_data = 12'heee;
			{8'd41, 8'd100}: color_data = 12'hbbb;
			{8'd41, 8'd101}: color_data = 12'heee;
			{8'd41, 8'd102}: color_data = 12'heee;
			{8'd41, 8'd103}: color_data = 12'hfff;
			{8'd41, 8'd104}: color_data = 12'hfff;
			{8'd41, 8'd105}: color_data = 12'heee;
			{8'd41, 8'd106}: color_data = 12'heee;
			{8'd41, 8'd107}: color_data = 12'h557;
			{8'd41, 8'd108}: color_data = 12'h249;
			{8'd41, 8'd109}: color_data = 12'h249;
			{8'd41, 8'd110}: color_data = 12'h249;
			{8'd41, 8'd111}: color_data = 12'h249;
			{8'd41, 8'd112}: color_data = 12'h247;
			{8'd41, 8'd113}: color_data = 12'h249;
			{8'd41, 8'd114}: color_data = 12'h249;
			{8'd41, 8'd115}: color_data = 12'h249;
			{8'd41, 8'd116}: color_data = 12'h249;
			{8'd41, 8'd117}: color_data = 12'h249;
			{8'd41, 8'd118}: color_data = 12'h249;
			{8'd41, 8'd119}: color_data = 12'h249;
			{8'd41, 8'd120}: color_data = 12'h248;
			{8'd41, 8'd121}: color_data = 12'h012;
			{8'd41, 8'd127}: color_data = 12'h000;
			{8'd41, 8'd128}: color_data = 12'h012;
			{8'd41, 8'd129}: color_data = 12'h024;
			{8'd41, 8'd130}: color_data = 12'h212;
			{8'd41, 8'd131}: color_data = 12'h532;
			{8'd41, 8'd132}: color_data = 12'h633;
			{8'd41, 8'd133}: color_data = 12'h643;
			{8'd41, 8'd134}: color_data = 12'h532;
			{8'd41, 8'd135}: color_data = 12'h643;
			{8'd41, 8'd136}: color_data = 12'h221;
			{8'd42, 8'd15}: color_data = 12'hfc5;
			{8'd42, 8'd16}: color_data = 12'hfc5;
			{8'd42, 8'd17}: color_data = 12'hfc4;
			{8'd42, 8'd18}: color_data = 12'hd90;
			{8'd42, 8'd19}: color_data = 12'hd90;
			{8'd42, 8'd20}: color_data = 12'hd90;
			{8'd42, 8'd21}: color_data = 12'hd90;
			{8'd42, 8'd22}: color_data = 12'hd90;
			{8'd42, 8'd23}: color_data = 12'hd90;
			{8'd42, 8'd24}: color_data = 12'hd90;
			{8'd42, 8'd25}: color_data = 12'hd90;
			{8'd42, 8'd26}: color_data = 12'hd90;
			{8'd42, 8'd27}: color_data = 12'hd90;
			{8'd42, 8'd28}: color_data = 12'hda0;
			{8'd42, 8'd29}: color_data = 12'hea1;
			{8'd42, 8'd30}: color_data = 12'heb3;
			{8'd42, 8'd31}: color_data = 12'hfc5;
			{8'd42, 8'd32}: color_data = 12'hfc5;
			{8'd42, 8'd33}: color_data = 12'hfc4;
			{8'd42, 8'd34}: color_data = 12'hff7;
			{8'd42, 8'd68}: color_data = 12'h110;
			{8'd42, 8'd69}: color_data = 12'h763;
			{8'd42, 8'd70}: color_data = 12'hb94;
			{8'd42, 8'd71}: color_data = 12'ha94;
			{8'd42, 8'd72}: color_data = 12'ha84;
			{8'd42, 8'd73}: color_data = 12'h864;
			{8'd42, 8'd74}: color_data = 12'hfdb;
			{8'd42, 8'd75}: color_data = 12'hfeb;
			{8'd42, 8'd76}: color_data = 12'hfdb;
			{8'd42, 8'd77}: color_data = 12'hfdb;
			{8'd42, 8'd78}: color_data = 12'hfdb;
			{8'd42, 8'd79}: color_data = 12'hfeb;
			{8'd42, 8'd80}: color_data = 12'hdb9;
			{8'd42, 8'd81}: color_data = 12'h455;
			{8'd42, 8'd82}: color_data = 12'h677;
			{8'd42, 8'd83}: color_data = 12'h566;
			{8'd42, 8'd84}: color_data = 12'h48a;
			{8'd42, 8'd85}: color_data = 12'h246;
			{8'd42, 8'd86}: color_data = 12'h001;
			{8'd42, 8'd87}: color_data = 12'h245;
			{8'd42, 8'd88}: color_data = 12'h49b;
			{8'd42, 8'd89}: color_data = 12'h48b;
			{8'd42, 8'd90}: color_data = 12'h378;
			{8'd42, 8'd91}: color_data = 12'h367;
			{8'd42, 8'd92}: color_data = 12'h357;
			{8'd42, 8'd93}: color_data = 12'h062;
			{8'd42, 8'd94}: color_data = 12'h0b3;
			{8'd42, 8'd95}: color_data = 12'h083;
			{8'd42, 8'd96}: color_data = 12'h586;
			{8'd42, 8'd97}: color_data = 12'h9aa;
			{8'd42, 8'd98}: color_data = 12'hbbb;
			{8'd42, 8'd99}: color_data = 12'haaa;
			{8'd42, 8'd100}: color_data = 12'haaa;
			{8'd42, 8'd101}: color_data = 12'haaa;
			{8'd42, 8'd102}: color_data = 12'haaa;
			{8'd42, 8'd103}: color_data = 12'hccc;
			{8'd42, 8'd104}: color_data = 12'hfff;
			{8'd42, 8'd105}: color_data = 12'hfff;
			{8'd42, 8'd106}: color_data = 12'hccc;
			{8'd42, 8'd107}: color_data = 12'h235;
			{8'd42, 8'd108}: color_data = 12'h248;
			{8'd42, 8'd109}: color_data = 12'h249;
			{8'd42, 8'd110}: color_data = 12'h249;
			{8'd42, 8'd111}: color_data = 12'h248;
			{8'd42, 8'd112}: color_data = 12'h136;
			{8'd42, 8'd113}: color_data = 12'h249;
			{8'd42, 8'd114}: color_data = 12'h249;
			{8'd42, 8'd115}: color_data = 12'h249;
			{8'd42, 8'd116}: color_data = 12'h249;
			{8'd42, 8'd117}: color_data = 12'h249;
			{8'd42, 8'd118}: color_data = 12'h249;
			{8'd42, 8'd119}: color_data = 12'h249;
			{8'd42, 8'd120}: color_data = 12'h249;
			{8'd42, 8'd121}: color_data = 12'h135;
			{8'd42, 8'd122}: color_data = 12'h000;
			{8'd42, 8'd125}: color_data = 12'h000;
			{8'd42, 8'd126}: color_data = 12'h012;
			{8'd42, 8'd127}: color_data = 12'h125;
			{8'd42, 8'd128}: color_data = 12'h248;
			{8'd42, 8'd129}: color_data = 12'h248;
			{8'd42, 8'd130}: color_data = 12'h422;
			{8'd42, 8'd131}: color_data = 12'h643;
			{8'd42, 8'd132}: color_data = 12'h633;
			{8'd42, 8'd133}: color_data = 12'h633;
			{8'd42, 8'd134}: color_data = 12'h643;
			{8'd42, 8'd135}: color_data = 12'hc96;
			{8'd42, 8'd136}: color_data = 12'h211;
			{8'd43, 8'd15}: color_data = 12'hfc5;
			{8'd43, 8'd16}: color_data = 12'hfc5;
			{8'd43, 8'd17}: color_data = 12'hfb3;
			{8'd43, 8'd18}: color_data = 12'hd90;
			{8'd43, 8'd19}: color_data = 12'hd90;
			{8'd43, 8'd20}: color_data = 12'hd90;
			{8'd43, 8'd21}: color_data = 12'hd90;
			{8'd43, 8'd22}: color_data = 12'hd90;
			{8'd43, 8'd23}: color_data = 12'hd90;
			{8'd43, 8'd24}: color_data = 12'hd90;
			{8'd43, 8'd25}: color_data = 12'hd90;
			{8'd43, 8'd26}: color_data = 12'hd90;
			{8'd43, 8'd27}: color_data = 12'hd90;
			{8'd43, 8'd28}: color_data = 12'hd90;
			{8'd43, 8'd29}: color_data = 12'hd90;
			{8'd43, 8'd30}: color_data = 12'hd90;
			{8'd43, 8'd31}: color_data = 12'hea1;
			{8'd43, 8'd32}: color_data = 12'hfc5;
			{8'd43, 8'd33}: color_data = 12'hfc5;
			{8'd43, 8'd34}: color_data = 12'hfd5;
			{8'd43, 8'd68}: color_data = 12'h210;
			{8'd43, 8'd69}: color_data = 12'hdb5;
			{8'd43, 8'd70}: color_data = 12'hfe7;
			{8'd43, 8'd71}: color_data = 12'hfe7;
			{8'd43, 8'd72}: color_data = 12'hfe7;
			{8'd43, 8'd73}: color_data = 12'ha84;
			{8'd43, 8'd74}: color_data = 12'h764;
			{8'd43, 8'd75}: color_data = 12'hba8;
			{8'd43, 8'd76}: color_data = 12'hdca;
			{8'd43, 8'd77}: color_data = 12'hfdb;
			{8'd43, 8'd78}: color_data = 12'heca;
			{8'd43, 8'd79}: color_data = 12'ha98;
			{8'd43, 8'd80}: color_data = 12'h467;
			{8'd43, 8'd81}: color_data = 12'h48a;
			{8'd43, 8'd82}: color_data = 12'h48a;
			{8'd43, 8'd83}: color_data = 12'h48a;
			{8'd43, 8'd84}: color_data = 12'h48a;
			{8'd43, 8'd85}: color_data = 12'h123;
			{8'd43, 8'd86}: color_data = 12'h001;
			{8'd43, 8'd87}: color_data = 12'h368;
			{8'd43, 8'd88}: color_data = 12'h49b;
			{8'd43, 8'd89}: color_data = 12'h48a;
			{8'd43, 8'd90}: color_data = 12'h48b;
			{8'd43, 8'd91}: color_data = 12'h367;
			{8'd43, 8'd92}: color_data = 12'h235;
			{8'd43, 8'd93}: color_data = 12'h144;
			{8'd43, 8'd94}: color_data = 12'h082;
			{8'd43, 8'd95}: color_data = 12'h0a3;
			{8'd43, 8'd96}: color_data = 12'h0a3;
			{8'd43, 8'd97}: color_data = 12'h062;
			{8'd43, 8'd98}: color_data = 12'hbaa;
			{8'd43, 8'd99}: color_data = 12'hfef;
			{8'd43, 8'd100}: color_data = 12'hfff;
			{8'd43, 8'd101}: color_data = 12'hfff;
			{8'd43, 8'd102}: color_data = 12'hfef;
			{8'd43, 8'd103}: color_data = 12'hede;
			{8'd43, 8'd104}: color_data = 12'hbcb;
			{8'd43, 8'd105}: color_data = 12'h797;
			{8'd43, 8'd106}: color_data = 12'h355;
			{8'd43, 8'd107}: color_data = 12'h368;
			{8'd43, 8'd108}: color_data = 12'h246;
			{8'd43, 8'd109}: color_data = 12'h136;
			{8'd43, 8'd110}: color_data = 12'h236;
			{8'd43, 8'd111}: color_data = 12'h124;
			{8'd43, 8'd112}: color_data = 12'h247;
			{8'd43, 8'd113}: color_data = 12'h249;
			{8'd43, 8'd114}: color_data = 12'h249;
			{8'd43, 8'd115}: color_data = 12'h249;
			{8'd43, 8'd116}: color_data = 12'h249;
			{8'd43, 8'd117}: color_data = 12'h249;
			{8'd43, 8'd118}: color_data = 12'h249;
			{8'd43, 8'd119}: color_data = 12'h249;
			{8'd43, 8'd120}: color_data = 12'h249;
			{8'd43, 8'd121}: color_data = 12'h248;
			{8'd43, 8'd122}: color_data = 12'h012;
			{8'd43, 8'd123}: color_data = 12'h000;
			{8'd43, 8'd124}: color_data = 12'h012;
			{8'd43, 8'd125}: color_data = 12'h135;
			{8'd43, 8'd126}: color_data = 12'h248;
			{8'd43, 8'd127}: color_data = 12'h249;
			{8'd43, 8'd128}: color_data = 12'h249;
			{8'd43, 8'd129}: color_data = 12'h136;
			{8'd43, 8'd130}: color_data = 12'h532;
			{8'd43, 8'd131}: color_data = 12'h643;
			{8'd43, 8'd132}: color_data = 12'h643;
			{8'd43, 8'd133}: color_data = 12'h532;
			{8'd43, 8'd134}: color_data = 12'ha85;
			{8'd43, 8'd135}: color_data = 12'ha85;
			{8'd43, 8'd136}: color_data = 12'h000;
			{8'd44, 8'd15}: color_data = 12'hfc5;
			{8'd44, 8'd16}: color_data = 12'hfc5;
			{8'd44, 8'd17}: color_data = 12'heb2;
			{8'd44, 8'd18}: color_data = 12'hd90;
			{8'd44, 8'd19}: color_data = 12'hd90;
			{8'd44, 8'd20}: color_data = 12'hd90;
			{8'd44, 8'd21}: color_data = 12'hd90;
			{8'd44, 8'd22}: color_data = 12'hd90;
			{8'd44, 8'd23}: color_data = 12'hd90;
			{8'd44, 8'd24}: color_data = 12'hd90;
			{8'd44, 8'd25}: color_data = 12'hd90;
			{8'd44, 8'd26}: color_data = 12'hd90;
			{8'd44, 8'd27}: color_data = 12'hd90;
			{8'd44, 8'd28}: color_data = 12'hd90;
			{8'd44, 8'd29}: color_data = 12'hd90;
			{8'd44, 8'd30}: color_data = 12'hd90;
			{8'd44, 8'd31}: color_data = 12'hea1;
			{8'd44, 8'd32}: color_data = 12'hfc5;
			{8'd44, 8'd33}: color_data = 12'hfc4;
			{8'd44, 8'd68}: color_data = 12'h331;
			{8'd44, 8'd69}: color_data = 12'h974;
			{8'd44, 8'd70}: color_data = 12'hb94;
			{8'd44, 8'd71}: color_data = 12'hca5;
			{8'd44, 8'd72}: color_data = 12'h984;
			{8'd44, 8'd73}: color_data = 12'hca5;
			{8'd44, 8'd74}: color_data = 12'hfd6;
			{8'd44, 8'd75}: color_data = 12'h873;
			{8'd44, 8'd76}: color_data = 12'hb95;
			{8'd44, 8'd77}: color_data = 12'h554;
			{8'd44, 8'd78}: color_data = 12'h367;
			{8'd44, 8'd79}: color_data = 12'h379;
			{8'd44, 8'd80}: color_data = 12'h48b;
			{8'd44, 8'd81}: color_data = 12'h48b;
			{8'd44, 8'd82}: color_data = 12'h48a;
			{8'd44, 8'd83}: color_data = 12'h48b;
			{8'd44, 8'd84}: color_data = 12'h479;
			{8'd44, 8'd85}: color_data = 12'h011;
			{8'd44, 8'd86}: color_data = 12'h012;
			{8'd44, 8'd87}: color_data = 12'h48a;
			{8'd44, 8'd88}: color_data = 12'h48b;
			{8'd44, 8'd89}: color_data = 12'h48a;
			{8'd44, 8'd90}: color_data = 12'h48a;
			{8'd44, 8'd91}: color_data = 12'h48b;
			{8'd44, 8'd92}: color_data = 12'h479;
			{8'd44, 8'd93}: color_data = 12'h47a;
			{8'd44, 8'd94}: color_data = 12'h255;
			{8'd44, 8'd95}: color_data = 12'h083;
			{8'd44, 8'd96}: color_data = 12'h0a3;
			{8'd44, 8'd97}: color_data = 12'h0a3;
			{8'd44, 8'd98}: color_data = 12'h174;
			{8'd44, 8'd99}: color_data = 12'h586;
			{8'd44, 8'd100}: color_data = 12'h687;
			{8'd44, 8'd101}: color_data = 12'h485;
			{8'd44, 8'd102}: color_data = 12'h274;
			{8'd44, 8'd103}: color_data = 12'h173;
			{8'd44, 8'd104}: color_data = 12'h082;
			{8'd44, 8'd105}: color_data = 12'h092;
			{8'd44, 8'd106}: color_data = 12'h164;
			{8'd44, 8'd107}: color_data = 12'h58b;
			{8'd44, 8'd108}: color_data = 12'h48b;
			{8'd44, 8'd109}: color_data = 12'h48a;
			{8'd44, 8'd110}: color_data = 12'h48a;
			{8'd44, 8'd111}: color_data = 12'h246;
			{8'd44, 8'd112}: color_data = 12'h248;
			{8'd44, 8'd113}: color_data = 12'h249;
			{8'd44, 8'd114}: color_data = 12'h249;
			{8'd44, 8'd115}: color_data = 12'h149;
			{8'd44, 8'd116}: color_data = 12'h149;
			{8'd44, 8'd117}: color_data = 12'h149;
			{8'd44, 8'd118}: color_data = 12'h149;
			{8'd44, 8'd119}: color_data = 12'h249;
			{8'd44, 8'd120}: color_data = 12'h249;
			{8'd44, 8'd121}: color_data = 12'h249;
			{8'd44, 8'd122}: color_data = 12'h137;
			{8'd44, 8'd123}: color_data = 12'h136;
			{8'd44, 8'd124}: color_data = 12'h248;
			{8'd44, 8'd125}: color_data = 12'h249;
			{8'd44, 8'd126}: color_data = 12'h249;
			{8'd44, 8'd127}: color_data = 12'h249;
			{8'd44, 8'd128}: color_data = 12'h249;
			{8'd44, 8'd129}: color_data = 12'h223;
			{8'd44, 8'd130}: color_data = 12'h633;
			{8'd44, 8'd131}: color_data = 12'h633;
			{8'd44, 8'd132}: color_data = 12'h633;
			{8'd44, 8'd133}: color_data = 12'h532;
			{8'd44, 8'd134}: color_data = 12'hda6;
			{8'd44, 8'd135}: color_data = 12'h974;
			{8'd44, 8'd136}: color_data = 12'h000;
			{8'd45, 8'd15}: color_data = 12'hfc4;
			{8'd45, 8'd16}: color_data = 12'hfc5;
			{8'd45, 8'd17}: color_data = 12'hea1;
			{8'd45, 8'd18}: color_data = 12'hd90;
			{8'd45, 8'd19}: color_data = 12'hd90;
			{8'd45, 8'd20}: color_data = 12'hd90;
			{8'd45, 8'd21}: color_data = 12'hea1;
			{8'd45, 8'd22}: color_data = 12'hfb3;
			{8'd45, 8'd23}: color_data = 12'hd90;
			{8'd45, 8'd24}: color_data = 12'hd90;
			{8'd45, 8'd25}: color_data = 12'hd90;
			{8'd45, 8'd26}: color_data = 12'hd90;
			{8'd45, 8'd27}: color_data = 12'hd90;
			{8'd45, 8'd28}: color_data = 12'hd90;
			{8'd45, 8'd29}: color_data = 12'hd90;
			{8'd45, 8'd30}: color_data = 12'hd90;
			{8'd45, 8'd31}: color_data = 12'heb2;
			{8'd45, 8'd32}: color_data = 12'hfc5;
			{8'd45, 8'd33}: color_data = 12'hfc4;
			{8'd45, 8'd68}: color_data = 12'h331;
			{8'd45, 8'd69}: color_data = 12'hba5;
			{8'd45, 8'd70}: color_data = 12'ha94;
			{8'd45, 8'd71}: color_data = 12'h652;
			{8'd45, 8'd72}: color_data = 12'hb94;
			{8'd45, 8'd73}: color_data = 12'hfe7;
			{8'd45, 8'd74}: color_data = 12'hfe7;
			{8'd45, 8'd75}: color_data = 12'ha84;
			{8'd45, 8'd76}: color_data = 12'ha94;
			{8'd45, 8'd77}: color_data = 12'h467;
			{8'd45, 8'd78}: color_data = 12'h49b;
			{8'd45, 8'd79}: color_data = 12'h48b;
			{8'd45, 8'd80}: color_data = 12'h48a;
			{8'd45, 8'd81}: color_data = 12'h48a;
			{8'd45, 8'd82}: color_data = 12'h48a;
			{8'd45, 8'd83}: color_data = 12'h49b;
			{8'd45, 8'd84}: color_data = 12'h256;
			{8'd45, 8'd85}: color_data = 12'h011;
			{8'd45, 8'd86}: color_data = 12'h012;
			{8'd45, 8'd87}: color_data = 12'h367;
			{8'd45, 8'd88}: color_data = 12'h49b;
			{8'd45, 8'd89}: color_data = 12'h48b;
			{8'd45, 8'd90}: color_data = 12'h48a;
			{8'd45, 8'd91}: color_data = 12'h48a;
			{8'd45, 8'd92}: color_data = 12'h48b;
			{8'd45, 8'd93}: color_data = 12'h48b;
			{8'd45, 8'd94}: color_data = 12'h48a;
			{8'd45, 8'd95}: color_data = 12'h154;
			{8'd45, 8'd96}: color_data = 12'h093;
			{8'd45, 8'd97}: color_data = 12'h0a3;
			{8'd45, 8'd98}: color_data = 12'h0a3;
			{8'd45, 8'd99}: color_data = 12'h0a3;
			{8'd45, 8'd100}: color_data = 12'h0a3;
			{8'd45, 8'd101}: color_data = 12'h0a3;
			{8'd45, 8'd102}: color_data = 12'h0a3;
			{8'd45, 8'd103}: color_data = 12'h0a3;
			{8'd45, 8'd104}: color_data = 12'h0a3;
			{8'd45, 8'd105}: color_data = 12'h0a3;
			{8'd45, 8'd106}: color_data = 12'h164;
			{8'd45, 8'd107}: color_data = 12'h48a;
			{8'd45, 8'd108}: color_data = 12'h48b;
			{8'd45, 8'd109}: color_data = 12'h48b;
			{8'd45, 8'd110}: color_data = 12'h59b;
			{8'd45, 8'd111}: color_data = 12'h257;
			{8'd45, 8'd112}: color_data = 12'h136;
			{8'd45, 8'd113}: color_data = 12'h236;
			{8'd45, 8'd114}: color_data = 12'h445;
			{8'd45, 8'd115}: color_data = 12'h655;
			{8'd45, 8'd116}: color_data = 12'h654;
			{8'd45, 8'd117}: color_data = 12'h654;
			{8'd45, 8'd118}: color_data = 12'h655;
			{8'd45, 8'd119}: color_data = 12'h445;
			{8'd45, 8'd120}: color_data = 12'h345;
			{8'd45, 8'd121}: color_data = 12'h236;
			{8'd45, 8'd122}: color_data = 12'h148;
			{8'd45, 8'd123}: color_data = 12'h149;
			{8'd45, 8'd124}: color_data = 12'h249;
			{8'd45, 8'd125}: color_data = 12'h249;
			{8'd45, 8'd126}: color_data = 12'h249;
			{8'd45, 8'd127}: color_data = 12'h249;
			{8'd45, 8'd128}: color_data = 12'h147;
			{8'd45, 8'd129}: color_data = 12'h422;
			{8'd45, 8'd130}: color_data = 12'h643;
			{8'd45, 8'd131}: color_data = 12'h633;
			{8'd45, 8'd132}: color_data = 12'h633;
			{8'd45, 8'd133}: color_data = 12'h643;
			{8'd45, 8'd134}: color_data = 12'heb7;
			{8'd45, 8'd135}: color_data = 12'h643;
			{8'd46, 8'd14}: color_data = 12'hcc6;
			{8'd46, 8'd15}: color_data = 12'hfc5;
			{8'd46, 8'd16}: color_data = 12'hfc5;
			{8'd46, 8'd17}: color_data = 12'hea1;
			{8'd46, 8'd18}: color_data = 12'hd90;
			{8'd46, 8'd19}: color_data = 12'hd90;
			{8'd46, 8'd20}: color_data = 12'hd90;
			{8'd46, 8'd21}: color_data = 12'heb3;
			{8'd46, 8'd22}: color_data = 12'hfc5;
			{8'd46, 8'd23}: color_data = 12'hd90;
			{8'd46, 8'd24}: color_data = 12'hd90;
			{8'd46, 8'd25}: color_data = 12'hd90;
			{8'd46, 8'd26}: color_data = 12'heb2;
			{8'd46, 8'd27}: color_data = 12'hea1;
			{8'd46, 8'd28}: color_data = 12'hd90;
			{8'd46, 8'd29}: color_data = 12'hd90;
			{8'd46, 8'd30}: color_data = 12'hd90;
			{8'd46, 8'd31}: color_data = 12'hfc4;
			{8'd46, 8'd32}: color_data = 12'hfc5;
			{8'd46, 8'd33}: color_data = 12'hfc5;
			{8'd46, 8'd67}: color_data = 12'h431;
			{8'd46, 8'd68}: color_data = 12'h763;
			{8'd46, 8'd69}: color_data = 12'h873;
			{8'd46, 8'd70}: color_data = 12'h653;
			{8'd46, 8'd71}: color_data = 12'h542;
			{8'd46, 8'd72}: color_data = 12'h652;
			{8'd46, 8'd73}: color_data = 12'ha84;
			{8'd46, 8'd74}: color_data = 12'ha94;
			{8'd46, 8'd75}: color_data = 12'h763;
			{8'd46, 8'd76}: color_data = 12'h344;
			{8'd46, 8'd77}: color_data = 12'h48b;
			{8'd46, 8'd78}: color_data = 12'h48b;
			{8'd46, 8'd79}: color_data = 12'h48a;
			{8'd46, 8'd80}: color_data = 12'h48a;
			{8'd46, 8'd81}: color_data = 12'h48a;
			{8'd46, 8'd82}: color_data = 12'h48a;
			{8'd46, 8'd83}: color_data = 12'h48b;
			{8'd46, 8'd84}: color_data = 12'h134;
			{8'd46, 8'd85}: color_data = 12'h001;
			{8'd46, 8'd86}: color_data = 12'h234;
			{8'd46, 8'd87}: color_data = 12'h368;
			{8'd46, 8'd88}: color_data = 12'h357;
			{8'd46, 8'd89}: color_data = 12'h48a;
			{8'd46, 8'd90}: color_data = 12'h48b;
			{8'd46, 8'd91}: color_data = 12'h48a;
			{8'd46, 8'd92}: color_data = 12'h48a;
			{8'd46, 8'd93}: color_data = 12'h48a;
			{8'd46, 8'd94}: color_data = 12'h48b;
			{8'd46, 8'd95}: color_data = 12'h48a;
			{8'd46, 8'd96}: color_data = 12'h154;
			{8'd46, 8'd97}: color_data = 12'h0a3;
			{8'd46, 8'd98}: color_data = 12'h0a3;
			{8'd46, 8'd99}: color_data = 12'h0a3;
			{8'd46, 8'd100}: color_data = 12'h0a3;
			{8'd46, 8'd101}: color_data = 12'h0a3;
			{8'd46, 8'd102}: color_data = 12'h0a3;
			{8'd46, 8'd103}: color_data = 12'h0a3;
			{8'd46, 8'd104}: color_data = 12'h0a3;
			{8'd46, 8'd105}: color_data = 12'h0a3;
			{8'd46, 8'd106}: color_data = 12'h164;
			{8'd46, 8'd107}: color_data = 12'h48a;
			{8'd46, 8'd108}: color_data = 12'h48a;
			{8'd46, 8'd109}: color_data = 12'h48b;
			{8'd46, 8'd110}: color_data = 12'h48a;
			{8'd46, 8'd111}: color_data = 12'h355;
			{8'd46, 8'd112}: color_data = 12'h964;
			{8'd46, 8'd113}: color_data = 12'hea5;
			{8'd46, 8'd114}: color_data = 12'hfb6;
			{8'd46, 8'd115}: color_data = 12'hfb6;
			{8'd46, 8'd116}: color_data = 12'hfb6;
			{8'd46, 8'd117}: color_data = 12'hfb6;
			{8'd46, 8'd118}: color_data = 12'hfb6;
			{8'd46, 8'd119}: color_data = 12'hfb6;
			{8'd46, 8'd120}: color_data = 12'hfa6;
			{8'd46, 8'd121}: color_data = 12'hd95;
			{8'd46, 8'd122}: color_data = 12'ha75;
			{8'd46, 8'd123}: color_data = 12'h654;
			{8'd46, 8'd124}: color_data = 12'h335;
			{8'd46, 8'd125}: color_data = 12'h148;
			{8'd46, 8'd126}: color_data = 12'h249;
			{8'd46, 8'd127}: color_data = 12'h249;
			{8'd46, 8'd128}: color_data = 12'h235;
			{8'd46, 8'd129}: color_data = 12'h532;
			{8'd46, 8'd130}: color_data = 12'h643;
			{8'd46, 8'd131}: color_data = 12'h643;
			{8'd46, 8'd132}: color_data = 12'h532;
			{8'd46, 8'd133}: color_data = 12'h864;
			{8'd46, 8'd134}: color_data = 12'hca6;
			{8'd46, 8'd135}: color_data = 12'h110;
			{8'd47, 8'd14}: color_data = 12'hfc4;
			{8'd47, 8'd15}: color_data = 12'hfc5;
			{8'd47, 8'd16}: color_data = 12'hfc4;
			{8'd47, 8'd17}: color_data = 12'hea0;
			{8'd47, 8'd18}: color_data = 12'hd90;
			{8'd47, 8'd19}: color_data = 12'hd90;
			{8'd47, 8'd20}: color_data = 12'hd90;
			{8'd47, 8'd21}: color_data = 12'hfc5;
			{8'd47, 8'd22}: color_data = 12'hfb4;
			{8'd47, 8'd23}: color_data = 12'hd90;
			{8'd47, 8'd24}: color_data = 12'hd90;
			{8'd47, 8'd25}: color_data = 12'hd90;
			{8'd47, 8'd26}: color_data = 12'hfc5;
			{8'd47, 8'd27}: color_data = 12'hea1;
			{8'd47, 8'd28}: color_data = 12'hd90;
			{8'd47, 8'd29}: color_data = 12'hd90;
			{8'd47, 8'd30}: color_data = 12'hd90;
			{8'd47, 8'd31}: color_data = 12'hfc4;
			{8'd47, 8'd32}: color_data = 12'hfc4;
			{8'd47, 8'd33}: color_data = 12'hfc5;
			{8'd47, 8'd66}: color_data = 12'h000;
			{8'd47, 8'd67}: color_data = 12'h763;
			{8'd47, 8'd68}: color_data = 12'h984;
			{8'd47, 8'd69}: color_data = 12'hb95;
			{8'd47, 8'd70}: color_data = 12'hec6;
			{8'd47, 8'd71}: color_data = 12'hdb5;
			{8'd47, 8'd72}: color_data = 12'h973;
			{8'd47, 8'd73}: color_data = 12'h763;
			{8'd47, 8'd74}: color_data = 12'ha84;
			{8'd47, 8'd75}: color_data = 12'h542;
			{8'd47, 8'd76}: color_data = 12'h378;
			{8'd47, 8'd77}: color_data = 12'h48b;
			{8'd47, 8'd78}: color_data = 12'h48a;
			{8'd47, 8'd79}: color_data = 12'h48a;
			{8'd47, 8'd80}: color_data = 12'h48a;
			{8'd47, 8'd81}: color_data = 12'h48a;
			{8'd47, 8'd82}: color_data = 12'h48b;
			{8'd47, 8'd83}: color_data = 12'h48a;
			{8'd47, 8'd84}: color_data = 12'h123;
			{8'd47, 8'd85}: color_data = 12'h011;
			{8'd47, 8'd86}: color_data = 12'h245;
			{8'd47, 8'd87}: color_data = 12'h59b;
			{8'd47, 8'd88}: color_data = 12'h479;
			{8'd47, 8'd89}: color_data = 12'h256;
			{8'd47, 8'd90}: color_data = 12'h368;
			{8'd47, 8'd91}: color_data = 12'h48a;
			{8'd47, 8'd92}: color_data = 12'h48a;
			{8'd47, 8'd93}: color_data = 12'h48a;
			{8'd47, 8'd94}: color_data = 12'h48a;
			{8'd47, 8'd95}: color_data = 12'h48b;
			{8'd47, 8'd96}: color_data = 12'h479;
			{8'd47, 8'd97}: color_data = 12'h063;
			{8'd47, 8'd98}: color_data = 12'h0a3;
			{8'd47, 8'd99}: color_data = 12'h0a3;
			{8'd47, 8'd100}: color_data = 12'h0a3;
			{8'd47, 8'd101}: color_data = 12'h0a3;
			{8'd47, 8'd102}: color_data = 12'h0a3;
			{8'd47, 8'd103}: color_data = 12'h0a3;
			{8'd47, 8'd104}: color_data = 12'h0a3;
			{8'd47, 8'd105}: color_data = 12'h0a3;
			{8'd47, 8'd106}: color_data = 12'h165;
			{8'd47, 8'd107}: color_data = 12'h48b;
			{8'd47, 8'd108}: color_data = 12'h48a;
			{8'd47, 8'd109}: color_data = 12'h48b;
			{8'd47, 8'd110}: color_data = 12'h456;
			{8'd47, 8'd111}: color_data = 12'hd95;
			{8'd47, 8'd112}: color_data = 12'hfb6;
			{8'd47, 8'd113}: color_data = 12'hfb6;
			{8'd47, 8'd114}: color_data = 12'hfb6;
			{8'd47, 8'd115}: color_data = 12'hfb6;
			{8'd47, 8'd116}: color_data = 12'hfb6;
			{8'd47, 8'd117}: color_data = 12'hfb6;
			{8'd47, 8'd118}: color_data = 12'hfb6;
			{8'd47, 8'd119}: color_data = 12'hfb6;
			{8'd47, 8'd120}: color_data = 12'hfb6;
			{8'd47, 8'd121}: color_data = 12'hfb6;
			{8'd47, 8'd122}: color_data = 12'hfb6;
			{8'd47, 8'd123}: color_data = 12'hfb6;
			{8'd47, 8'd124}: color_data = 12'hea5;
			{8'd47, 8'd125}: color_data = 12'h864;
			{8'd47, 8'd126}: color_data = 12'h236;
			{8'd47, 8'd127}: color_data = 12'h148;
			{8'd47, 8'd128}: color_data = 12'h323;
			{8'd47, 8'd129}: color_data = 12'h633;
			{8'd47, 8'd130}: color_data = 12'h633;
			{8'd47, 8'd131}: color_data = 12'h643;
			{8'd47, 8'd132}: color_data = 12'h422;
			{8'd47, 8'd133}: color_data = 12'h221;
			{8'd47, 8'd134}: color_data = 12'h864;
			{8'd47, 8'd135}: color_data = 12'h110;
			{8'd48, 8'd14}: color_data = 12'hfc4;
			{8'd48, 8'd15}: color_data = 12'hfc4;
			{8'd48, 8'd16}: color_data = 12'hfb3;
			{8'd48, 8'd17}: color_data = 12'hd90;
			{8'd48, 8'd18}: color_data = 12'hd90;
			{8'd48, 8'd19}: color_data = 12'hd90;
			{8'd48, 8'd20}: color_data = 12'hea1;
			{8'd48, 8'd21}: color_data = 12'hfc6;
			{8'd48, 8'd22}: color_data = 12'hfb3;
			{8'd48, 8'd23}: color_data = 12'hd90;
			{8'd48, 8'd24}: color_data = 12'hd90;
			{8'd48, 8'd25}: color_data = 12'hea1;
			{8'd48, 8'd26}: color_data = 12'hfc5;
			{8'd48, 8'd27}: color_data = 12'hea0;
			{8'd48, 8'd28}: color_data = 12'hd90;
			{8'd48, 8'd29}: color_data = 12'hd90;
			{8'd48, 8'd30}: color_data = 12'hea1;
			{8'd48, 8'd31}: color_data = 12'hfc5;
			{8'd48, 8'd32}: color_data = 12'hfc5;
			{8'd48, 8'd33}: color_data = 12'hfb7;
			{8'd48, 8'd66}: color_data = 12'h000;
			{8'd48, 8'd67}: color_data = 12'h652;
			{8'd48, 8'd68}: color_data = 12'hdb5;
			{8'd48, 8'd69}: color_data = 12'hfe7;
			{8'd48, 8'd70}: color_data = 12'hfd7;
			{8'd48, 8'd71}: color_data = 12'hfe7;
			{8'd48, 8'd72}: color_data = 12'hba5;
			{8'd48, 8'd73}: color_data = 12'h984;
			{8'd48, 8'd74}: color_data = 12'hdb5;
			{8'd48, 8'd75}: color_data = 12'h775;
			{8'd48, 8'd76}: color_data = 12'h48a;
			{8'd48, 8'd77}: color_data = 12'h48b;
			{8'd48, 8'd78}: color_data = 12'h48a;
			{8'd48, 8'd79}: color_data = 12'h48a;
			{8'd48, 8'd80}: color_data = 12'h48a;
			{8'd48, 8'd81}: color_data = 12'h48a;
			{8'd48, 8'd82}: color_data = 12'h48b;
			{8'd48, 8'd83}: color_data = 12'h48a;
			{8'd48, 8'd84}: color_data = 12'h112;
			{8'd48, 8'd85}: color_data = 12'h011;
			{8'd48, 8'd86}: color_data = 12'h357;
			{8'd48, 8'd87}: color_data = 12'h49b;
			{8'd48, 8'd88}: color_data = 12'h48b;
			{8'd48, 8'd89}: color_data = 12'h48b;
			{8'd48, 8'd90}: color_data = 12'h48a;
			{8'd48, 8'd91}: color_data = 12'h48a;
			{8'd48, 8'd92}: color_data = 12'h48a;
			{8'd48, 8'd93}: color_data = 12'h48a;
			{8'd48, 8'd94}: color_data = 12'h48a;
			{8'd48, 8'd95}: color_data = 12'h48a;
			{8'd48, 8'd96}: color_data = 12'h49b;
			{8'd48, 8'd97}: color_data = 12'h368;
			{8'd48, 8'd98}: color_data = 12'h063;
			{8'd48, 8'd99}: color_data = 12'h0a3;
			{8'd48, 8'd100}: color_data = 12'h0a3;
			{8'd48, 8'd101}: color_data = 12'h0a3;
			{8'd48, 8'd102}: color_data = 12'h0a3;
			{8'd48, 8'd103}: color_data = 12'h0a3;
			{8'd48, 8'd104}: color_data = 12'h0a3;
			{8'd48, 8'd105}: color_data = 12'h083;
			{8'd48, 8'd106}: color_data = 12'h367;
			{8'd48, 8'd107}: color_data = 12'h48b;
			{8'd48, 8'd108}: color_data = 12'h48b;
			{8'd48, 8'd109}: color_data = 12'h368;
			{8'd48, 8'd110}: color_data = 12'hb84;
			{8'd48, 8'd111}: color_data = 12'hfb6;
			{8'd48, 8'd112}: color_data = 12'hfb6;
			{8'd48, 8'd113}: color_data = 12'hfb6;
			{8'd48, 8'd114}: color_data = 12'hfb6;
			{8'd48, 8'd115}: color_data = 12'hfb6;
			{8'd48, 8'd116}: color_data = 12'hfb6;
			{8'd48, 8'd117}: color_data = 12'hfb6;
			{8'd48, 8'd118}: color_data = 12'hfb6;
			{8'd48, 8'd119}: color_data = 12'hfb6;
			{8'd48, 8'd120}: color_data = 12'hfb6;
			{8'd48, 8'd121}: color_data = 12'hfb6;
			{8'd48, 8'd122}: color_data = 12'hfb6;
			{8'd48, 8'd123}: color_data = 12'hfb6;
			{8'd48, 8'd124}: color_data = 12'hfb6;
			{8'd48, 8'd125}: color_data = 12'hfb6;
			{8'd48, 8'd126}: color_data = 12'hc95;
			{8'd48, 8'd127}: color_data = 12'h334;
			{8'd48, 8'd128}: color_data = 12'h422;
			{8'd48, 8'd129}: color_data = 12'h643;
			{8'd48, 8'd130}: color_data = 12'h633;
			{8'd48, 8'd131}: color_data = 12'h533;
			{8'd48, 8'd132}: color_data = 12'h643;
			{8'd48, 8'd133}: color_data = 12'h874;
			{8'd48, 8'd134}: color_data = 12'h000;
			{8'd49, 8'd14}: color_data = 12'hfc5;
			{8'd49, 8'd15}: color_data = 12'hfc4;
			{8'd49, 8'd16}: color_data = 12'hfc4;
			{8'd49, 8'd17}: color_data = 12'hfc3;
			{8'd49, 8'd18}: color_data = 12'hfb3;
			{8'd49, 8'd19}: color_data = 12'hfb3;
			{8'd49, 8'd20}: color_data = 12'hfc4;
			{8'd49, 8'd21}: color_data = 12'hfc5;
			{8'd49, 8'd22}: color_data = 12'hfc5;
			{8'd49, 8'd23}: color_data = 12'hfc4;
			{8'd49, 8'd24}: color_data = 12'hfb3;
			{8'd49, 8'd25}: color_data = 12'hfc4;
			{8'd49, 8'd26}: color_data = 12'hfc4;
			{8'd49, 8'd27}: color_data = 12'hd90;
			{8'd49, 8'd28}: color_data = 12'hd90;
			{8'd49, 8'd29}: color_data = 12'hd90;
			{8'd49, 8'd30}: color_data = 12'hea2;
			{8'd49, 8'd31}: color_data = 12'hfc5;
			{8'd49, 8'd32}: color_data = 12'hfc5;
			{8'd49, 8'd67}: color_data = 12'h321;
			{8'd49, 8'd68}: color_data = 12'hcb5;
			{8'd49, 8'd69}: color_data = 12'hfd7;
			{8'd49, 8'd70}: color_data = 12'hfd6;
			{8'd49, 8'd71}: color_data = 12'hca5;
			{8'd49, 8'd72}: color_data = 12'h984;
			{8'd49, 8'd73}: color_data = 12'hfe7;
			{8'd49, 8'd74}: color_data = 12'hfd6;
			{8'd49, 8'd75}: color_data = 12'h566;
			{8'd49, 8'd76}: color_data = 12'h48b;
			{8'd49, 8'd77}: color_data = 12'h48a;
			{8'd49, 8'd78}: color_data = 12'h48a;
			{8'd49, 8'd79}: color_data = 12'h48a;
			{8'd49, 8'd80}: color_data = 12'h48a;
			{8'd49, 8'd81}: color_data = 12'h48a;
			{8'd49, 8'd82}: color_data = 12'h48b;
			{8'd49, 8'd83}: color_data = 12'h479;
			{8'd49, 8'd84}: color_data = 12'h112;
			{8'd49, 8'd85}: color_data = 12'h011;
			{8'd49, 8'd86}: color_data = 12'h245;
			{8'd49, 8'd87}: color_data = 12'h48b;
			{8'd49, 8'd88}: color_data = 12'h48b;
			{8'd49, 8'd89}: color_data = 12'h48a;
			{8'd49, 8'd90}: color_data = 12'h48b;
			{8'd49, 8'd91}: color_data = 12'h48a;
			{8'd49, 8'd92}: color_data = 12'h48a;
			{8'd49, 8'd93}: color_data = 12'h48a;
			{8'd49, 8'd94}: color_data = 12'h48a;
			{8'd49, 8'd95}: color_data = 12'h48a;
			{8'd49, 8'd96}: color_data = 12'h48a;
			{8'd49, 8'd97}: color_data = 12'h49b;
			{8'd49, 8'd98}: color_data = 12'h368;
			{8'd49, 8'd99}: color_data = 12'h072;
			{8'd49, 8'd100}: color_data = 12'h0a3;
			{8'd49, 8'd101}: color_data = 12'h0a3;
			{8'd49, 8'd102}: color_data = 12'h0a3;
			{8'd49, 8'd103}: color_data = 12'h0a3;
			{8'd49, 8'd104}: color_data = 12'h0a3;
			{8'd49, 8'd105}: color_data = 12'h063;
			{8'd49, 8'd106}: color_data = 12'h47a;
			{8'd49, 8'd107}: color_data = 12'h48b;
			{8'd49, 8'd108}: color_data = 12'h48a;
			{8'd49, 8'd109}: color_data = 12'h665;
			{8'd49, 8'd110}: color_data = 12'hfb6;
			{8'd49, 8'd111}: color_data = 12'hfb6;
			{8'd49, 8'd112}: color_data = 12'hfb6;
			{8'd49, 8'd113}: color_data = 12'hfb6;
			{8'd49, 8'd114}: color_data = 12'hfb6;
			{8'd49, 8'd115}: color_data = 12'hfb6;
			{8'd49, 8'd116}: color_data = 12'hfb6;
			{8'd49, 8'd117}: color_data = 12'hfb6;
			{8'd49, 8'd118}: color_data = 12'hfb6;
			{8'd49, 8'd119}: color_data = 12'hfb6;
			{8'd49, 8'd120}: color_data = 12'hfb6;
			{8'd49, 8'd121}: color_data = 12'hfb6;
			{8'd49, 8'd122}: color_data = 12'hfb6;
			{8'd49, 8'd123}: color_data = 12'hfb6;
			{8'd49, 8'd124}: color_data = 12'hfb6;
			{8'd49, 8'd125}: color_data = 12'hfb6;
			{8'd49, 8'd126}: color_data = 12'hfb6;
			{8'd49, 8'd127}: color_data = 12'hd95;
			{8'd49, 8'd128}: color_data = 12'h532;
			{8'd49, 8'd129}: color_data = 12'h633;
			{8'd49, 8'd130}: color_data = 12'h643;
			{8'd49, 8'd131}: color_data = 12'h432;
			{8'd49, 8'd132}: color_data = 12'hb95;
			{8'd49, 8'd133}: color_data = 12'hb95;
			{8'd49, 8'd134}: color_data = 12'h110;
			{8'd50, 8'd14}: color_data = 12'hf77;
			{8'd50, 8'd15}: color_data = 12'hfc4;
			{8'd50, 8'd16}: color_data = 12'hfc5;
			{8'd50, 8'd17}: color_data = 12'hfc5;
			{8'd50, 8'd18}: color_data = 12'hfc5;
			{8'd50, 8'd19}: color_data = 12'hfc5;
			{8'd50, 8'd20}: color_data = 12'hfc5;
			{8'd50, 8'd21}: color_data = 12'hfc5;
			{8'd50, 8'd22}: color_data = 12'hfc4;
			{8'd50, 8'd23}: color_data = 12'hfc5;
			{8'd50, 8'd24}: color_data = 12'hfc6;
			{8'd50, 8'd25}: color_data = 12'hfc6;
			{8'd50, 8'd26}: color_data = 12'hfb4;
			{8'd50, 8'd27}: color_data = 12'hd90;
			{8'd50, 8'd28}: color_data = 12'hd90;
			{8'd50, 8'd29}: color_data = 12'hd90;
			{8'd50, 8'd30}: color_data = 12'heb3;
			{8'd50, 8'd31}: color_data = 12'hfc5;
			{8'd50, 8'd32}: color_data = 12'hfc5;
			{8'd50, 8'd67}: color_data = 12'h000;
			{8'd50, 8'd68}: color_data = 12'h221;
			{8'd50, 8'd69}: color_data = 12'h652;
			{8'd50, 8'd70}: color_data = 12'h542;
			{8'd50, 8'd71}: color_data = 12'h000;
			{8'd50, 8'd72}: color_data = 12'h552;
			{8'd50, 8'd73}: color_data = 12'h984;
			{8'd50, 8'd74}: color_data = 12'h652;
			{8'd50, 8'd75}: color_data = 12'h367;
			{8'd50, 8'd76}: color_data = 12'h49b;
			{8'd50, 8'd77}: color_data = 12'h48a;
			{8'd50, 8'd78}: color_data = 12'h48b;
			{8'd50, 8'd79}: color_data = 12'h48a;
			{8'd50, 8'd80}: color_data = 12'h48a;
			{8'd50, 8'd81}: color_data = 12'h48a;
			{8'd50, 8'd82}: color_data = 12'h48b;
			{8'd50, 8'd83}: color_data = 12'h48a;
			{8'd50, 8'd84}: color_data = 12'h112;
			{8'd50, 8'd85}: color_data = 12'h011;
			{8'd50, 8'd86}: color_data = 12'h246;
			{8'd50, 8'd87}: color_data = 12'h357;
			{8'd50, 8'd88}: color_data = 12'h48a;
			{8'd50, 8'd89}: color_data = 12'h48b;
			{8'd50, 8'd90}: color_data = 12'h48a;
			{8'd50, 8'd91}: color_data = 12'h48a;
			{8'd50, 8'd92}: color_data = 12'h48a;
			{8'd50, 8'd93}: color_data = 12'h48a;
			{8'd50, 8'd94}: color_data = 12'h48a;
			{8'd50, 8'd95}: color_data = 12'h48a;
			{8'd50, 8'd96}: color_data = 12'h48a;
			{8'd50, 8'd97}: color_data = 12'h48a;
			{8'd50, 8'd98}: color_data = 12'h48b;
			{8'd50, 8'd99}: color_data = 12'h367;
			{8'd50, 8'd100}: color_data = 12'h072;
			{8'd50, 8'd101}: color_data = 12'h0a3;
			{8'd50, 8'd102}: color_data = 12'h0a3;
			{8'd50, 8'd103}: color_data = 12'h0a3;
			{8'd50, 8'd104}: color_data = 12'h082;
			{8'd50, 8'd105}: color_data = 12'h266;
			{8'd50, 8'd106}: color_data = 12'h48b;
			{8'd50, 8'd107}: color_data = 12'h48b;
			{8'd50, 8'd108}: color_data = 12'h48a;
			{8'd50, 8'd109}: color_data = 12'h443;
			{8'd50, 8'd110}: color_data = 12'hea5;
			{8'd50, 8'd111}: color_data = 12'hfb6;
			{8'd50, 8'd112}: color_data = 12'hfb6;
			{8'd50, 8'd113}: color_data = 12'hfb6;
			{8'd50, 8'd114}: color_data = 12'hfb6;
			{8'd50, 8'd115}: color_data = 12'hfb6;
			{8'd50, 8'd116}: color_data = 12'hfb6;
			{8'd50, 8'd117}: color_data = 12'hfb6;
			{8'd50, 8'd118}: color_data = 12'hfb6;
			{8'd50, 8'd119}: color_data = 12'hfb6;
			{8'd50, 8'd120}: color_data = 12'hfb6;
			{8'd50, 8'd121}: color_data = 12'hfb6;
			{8'd50, 8'd122}: color_data = 12'hfb6;
			{8'd50, 8'd123}: color_data = 12'hfb6;
			{8'd50, 8'd124}: color_data = 12'hfb6;
			{8'd50, 8'd125}: color_data = 12'hfb6;
			{8'd50, 8'd126}: color_data = 12'hfb6;
			{8'd50, 8'd127}: color_data = 12'hfb6;
			{8'd50, 8'd128}: color_data = 12'hb84;
			{8'd50, 8'd129}: color_data = 12'h432;
			{8'd50, 8'd130}: color_data = 12'h533;
			{8'd50, 8'd131}: color_data = 12'h653;
			{8'd50, 8'd132}: color_data = 12'heb7;
			{8'd50, 8'd133}: color_data = 12'h864;
			{8'd50, 8'd134}: color_data = 12'h000;
			{8'd51, 8'd15}: color_data = 12'hff7;
			{8'd51, 8'd16}: color_data = 12'hfc5;
			{8'd51, 8'd17}: color_data = 12'hfc5;
			{8'd51, 8'd18}: color_data = 12'hfc6;
			{8'd51, 8'd19}: color_data = 12'hfc5;
			{8'd51, 8'd20}: color_data = 12'hfc5;
			{8'd51, 8'd21}: color_data = 12'hfc6;
			{8'd51, 8'd22}: color_data = 12'hfc6;
			{8'd51, 8'd23}: color_data = 12'hfc5;
			{8'd51, 8'd24}: color_data = 12'hfc5;
			{8'd51, 8'd25}: color_data = 12'hfc4;
			{8'd51, 8'd26}: color_data = 12'hfc4;
			{8'd51, 8'd27}: color_data = 12'hfb2;
			{8'd51, 8'd28}: color_data = 12'hd90;
			{8'd51, 8'd29}: color_data = 12'hd90;
			{8'd51, 8'd30}: color_data = 12'hfc4;
			{8'd51, 8'd31}: color_data = 12'hfc5;
			{8'd51, 8'd32}: color_data = 12'hfc4;
			{8'd51, 8'd74}: color_data = 12'h000;
			{8'd51, 8'd75}: color_data = 12'h368;
			{8'd51, 8'd76}: color_data = 12'h59b;
			{8'd51, 8'd77}: color_data = 12'h49b;
			{8'd51, 8'd78}: color_data = 12'h48a;
			{8'd51, 8'd79}: color_data = 12'h48a;
			{8'd51, 8'd80}: color_data = 12'h48a;
			{8'd51, 8'd81}: color_data = 12'h48a;
			{8'd51, 8'd82}: color_data = 12'h49b;
			{8'd51, 8'd83}: color_data = 12'h479;
			{8'd51, 8'd84}: color_data = 12'h012;
			{8'd51, 8'd85}: color_data = 12'h011;
			{8'd51, 8'd86}: color_data = 12'h368;
			{8'd51, 8'd87}: color_data = 12'h479;
			{8'd51, 8'd88}: color_data = 12'h256;
			{8'd51, 8'd89}: color_data = 12'h479;
			{8'd51, 8'd90}: color_data = 12'h48b;
			{8'd51, 8'd91}: color_data = 12'h48a;
			{8'd51, 8'd92}: color_data = 12'h48a;
			{8'd51, 8'd93}: color_data = 12'h48a;
			{8'd51, 8'd94}: color_data = 12'h48a;
			{8'd51, 8'd95}: color_data = 12'h48a;
			{8'd51, 8'd96}: color_data = 12'h48a;
			{8'd51, 8'd97}: color_data = 12'h48a;
			{8'd51, 8'd98}: color_data = 12'h48a;
			{8'd51, 8'd99}: color_data = 12'h48b;
			{8'd51, 8'd100}: color_data = 12'h368;
			{8'd51, 8'd101}: color_data = 12'h164;
			{8'd51, 8'd102}: color_data = 12'h082;
			{8'd51, 8'd103}: color_data = 12'h073;
			{8'd51, 8'd104}: color_data = 12'h256;
			{8'd51, 8'd105}: color_data = 12'h48a;
			{8'd51, 8'd106}: color_data = 12'h48b;
			{8'd51, 8'd107}: color_data = 12'h48a;
			{8'd51, 8'd108}: color_data = 12'h48b;
			{8'd51, 8'd109}: color_data = 12'h333;
			{8'd51, 8'd110}: color_data = 12'h632;
			{8'd51, 8'd111}: color_data = 12'hc95;
			{8'd51, 8'd112}: color_data = 12'hfb6;
			{8'd51, 8'd113}: color_data = 12'hfb6;
			{8'd51, 8'd114}: color_data = 12'hfb6;
			{8'd51, 8'd115}: color_data = 12'hfb6;
			{8'd51, 8'd116}: color_data = 12'hfb6;
			{8'd51, 8'd117}: color_data = 12'hfb6;
			{8'd51, 8'd118}: color_data = 12'hfb6;
			{8'd51, 8'd119}: color_data = 12'hfb6;
			{8'd51, 8'd120}: color_data = 12'hfb6;
			{8'd51, 8'd121}: color_data = 12'hfb6;
			{8'd51, 8'd122}: color_data = 12'hfb6;
			{8'd51, 8'd123}: color_data = 12'hfb6;
			{8'd51, 8'd124}: color_data = 12'hfb6;
			{8'd51, 8'd125}: color_data = 12'hfb6;
			{8'd51, 8'd126}: color_data = 12'hfb6;
			{8'd51, 8'd127}: color_data = 12'hfb6;
			{8'd51, 8'd128}: color_data = 12'hfb6;
			{8'd51, 8'd129}: color_data = 12'h753;
			{8'd51, 8'd130}: color_data = 12'h321;
			{8'd51, 8'd131}: color_data = 12'hb95;
			{8'd51, 8'd132}: color_data = 12'heb7;
			{8'd51, 8'd133}: color_data = 12'h542;
			{8'd52, 8'd25}: color_data = 12'hfc4;
			{8'd52, 8'd26}: color_data = 12'hfc4;
			{8'd52, 8'd27}: color_data = 12'hfc5;
			{8'd52, 8'd28}: color_data = 12'hfb3;
			{8'd52, 8'd29}: color_data = 12'hea1;
			{8'd52, 8'd30}: color_data = 12'hfc5;
			{8'd52, 8'd31}: color_data = 12'hfc5;
			{8'd52, 8'd32}: color_data = 12'hfc4;
			{8'd52, 8'd74}: color_data = 12'h000;
			{8'd52, 8'd75}: color_data = 12'h134;
			{8'd52, 8'd76}: color_data = 12'h356;
			{8'd52, 8'd77}: color_data = 12'h245;
			{8'd52, 8'd78}: color_data = 12'h112;
			{8'd52, 8'd79}: color_data = 12'h367;
			{8'd52, 8'd80}: color_data = 12'h59b;
			{8'd52, 8'd81}: color_data = 12'h49b;
			{8'd52, 8'd82}: color_data = 12'h368;
			{8'd52, 8'd83}: color_data = 12'h112;
			{8'd52, 8'd84}: color_data = 12'h001;
			{8'd52, 8'd85}: color_data = 12'h011;
			{8'd52, 8'd86}: color_data = 12'h368;
			{8'd52, 8'd87}: color_data = 12'h49b;
			{8'd52, 8'd88}: color_data = 12'h48a;
			{8'd52, 8'd89}: color_data = 12'h48a;
			{8'd52, 8'd90}: color_data = 12'h48b;
			{8'd52, 8'd91}: color_data = 12'h48a;
			{8'd52, 8'd92}: color_data = 12'h48a;
			{8'd52, 8'd93}: color_data = 12'h48a;
			{8'd52, 8'd94}: color_data = 12'h48a;
			{8'd52, 8'd95}: color_data = 12'h48a;
			{8'd52, 8'd96}: color_data = 12'h48a;
			{8'd52, 8'd97}: color_data = 12'h48a;
			{8'd52, 8'd98}: color_data = 12'h48a;
			{8'd52, 8'd99}: color_data = 12'h48a;
			{8'd52, 8'd100}: color_data = 12'h48b;
			{8'd52, 8'd101}: color_data = 12'h48a;
			{8'd52, 8'd102}: color_data = 12'h378;
			{8'd52, 8'd103}: color_data = 12'h479;
			{8'd52, 8'd104}: color_data = 12'h48b;
			{8'd52, 8'd105}: color_data = 12'h48b;
			{8'd52, 8'd106}: color_data = 12'h48a;
			{8'd52, 8'd107}: color_data = 12'h48a;
			{8'd52, 8'd108}: color_data = 12'h49b;
			{8'd52, 8'd109}: color_data = 12'h356;
			{8'd52, 8'd110}: color_data = 12'h732;
			{8'd52, 8'd111}: color_data = 12'h632;
			{8'd52, 8'd112}: color_data = 12'hb74;
			{8'd52, 8'd113}: color_data = 12'hfb6;
			{8'd52, 8'd114}: color_data = 12'hfb6;
			{8'd52, 8'd115}: color_data = 12'hfb6;
			{8'd52, 8'd116}: color_data = 12'hfb6;
			{8'd52, 8'd117}: color_data = 12'hfb6;
			{8'd52, 8'd118}: color_data = 12'hfb6;
			{8'd52, 8'd119}: color_data = 12'hfb6;
			{8'd52, 8'd120}: color_data = 12'hfb6;
			{8'd52, 8'd121}: color_data = 12'hfb6;
			{8'd52, 8'd122}: color_data = 12'hfb6;
			{8'd52, 8'd123}: color_data = 12'hfb6;
			{8'd52, 8'd124}: color_data = 12'hfb6;
			{8'd52, 8'd125}: color_data = 12'hfb6;
			{8'd52, 8'd126}: color_data = 12'hfb6;
			{8'd52, 8'd127}: color_data = 12'hfb6;
			{8'd52, 8'd128}: color_data = 12'hfb6;
			{8'd52, 8'd129}: color_data = 12'ha74;
			{8'd52, 8'd130}: color_data = 12'h963;
			{8'd52, 8'd131}: color_data = 12'h753;
			{8'd52, 8'd132}: color_data = 12'h974;
			{8'd52, 8'd133}: color_data = 12'h211;
			{8'd53, 8'd26}: color_data = 12'hfc4;
			{8'd53, 8'd27}: color_data = 12'hfc4;
			{8'd53, 8'd28}: color_data = 12'hfc5;
			{8'd53, 8'd29}: color_data = 12'hfc5;
			{8'd53, 8'd30}: color_data = 12'hfc5;
			{8'd53, 8'd31}: color_data = 12'hfc5;
			{8'd53, 8'd75}: color_data = 12'h000;
			{8'd53, 8'd76}: color_data = 12'h000;
			{8'd53, 8'd77}: color_data = 12'h000;
			{8'd53, 8'd79}: color_data = 12'h122;
			{8'd53, 8'd80}: color_data = 12'h367;
			{8'd53, 8'd81}: color_data = 12'h256;
			{8'd53, 8'd82}: color_data = 12'h011;
			{8'd53, 8'd84}: color_data = 12'h000;
			{8'd53, 8'd85}: color_data = 12'h000;
			{8'd53, 8'd86}: color_data = 12'h367;
			{8'd53, 8'd87}: color_data = 12'h59b;
			{8'd53, 8'd88}: color_data = 12'h48a;
			{8'd53, 8'd89}: color_data = 12'h48b;
			{8'd53, 8'd90}: color_data = 12'h48a;
			{8'd53, 8'd91}: color_data = 12'h48a;
			{8'd53, 8'd92}: color_data = 12'h48a;
			{8'd53, 8'd93}: color_data = 12'h48a;
			{8'd53, 8'd94}: color_data = 12'h48a;
			{8'd53, 8'd95}: color_data = 12'h48a;
			{8'd53, 8'd96}: color_data = 12'h48a;
			{8'd53, 8'd97}: color_data = 12'h48a;
			{8'd53, 8'd98}: color_data = 12'h48a;
			{8'd53, 8'd99}: color_data = 12'h48a;
			{8'd53, 8'd100}: color_data = 12'h48a;
			{8'd53, 8'd101}: color_data = 12'h48b;
			{8'd53, 8'd102}: color_data = 12'h48b;
			{8'd53, 8'd103}: color_data = 12'h48b;
			{8'd53, 8'd104}: color_data = 12'h48a;
			{8'd53, 8'd105}: color_data = 12'h48a;
			{8'd53, 8'd106}: color_data = 12'h48a;
			{8'd53, 8'd107}: color_data = 12'h48a;
			{8'd53, 8'd108}: color_data = 12'h48b;
			{8'd53, 8'd109}: color_data = 12'h479;
			{8'd53, 8'd110}: color_data = 12'h532;
			{8'd53, 8'd111}: color_data = 12'h842;
			{8'd53, 8'd112}: color_data = 12'h632;
			{8'd53, 8'd113}: color_data = 12'h963;
			{8'd53, 8'd114}: color_data = 12'hfb6;
			{8'd53, 8'd115}: color_data = 12'hfb6;
			{8'd53, 8'd116}: color_data = 12'hfb6;
			{8'd53, 8'd117}: color_data = 12'hfb6;
			{8'd53, 8'd118}: color_data = 12'hfb6;
			{8'd53, 8'd119}: color_data = 12'hfb6;
			{8'd53, 8'd120}: color_data = 12'hfb6;
			{8'd53, 8'd121}: color_data = 12'hfb6;
			{8'd53, 8'd122}: color_data = 12'hfb6;
			{8'd53, 8'd123}: color_data = 12'hfb6;
			{8'd53, 8'd124}: color_data = 12'hfb6;
			{8'd53, 8'd125}: color_data = 12'hfb6;
			{8'd53, 8'd126}: color_data = 12'hfb6;
			{8'd53, 8'd127}: color_data = 12'hfb6;
			{8'd53, 8'd128}: color_data = 12'hfb6;
			{8'd53, 8'd129}: color_data = 12'ha74;
			{8'd53, 8'd130}: color_data = 12'hc95;
			{8'd53, 8'd131}: color_data = 12'hb84;
			{8'd53, 8'd132}: color_data = 12'hd95;
			{8'd53, 8'd133}: color_data = 12'h753;
			{8'd53, 8'd134}: color_data = 12'h000;
			{8'd54, 8'd27}: color_data = 12'hfc6;
			{8'd54, 8'd28}: color_data = 12'hfc4;
			{8'd54, 8'd29}: color_data = 12'hfc5;
			{8'd54, 8'd30}: color_data = 12'hfc5;
			{8'd54, 8'd31}: color_data = 12'hfc5;
			{8'd54, 8'd79}: color_data = 12'h000;
			{8'd54, 8'd80}: color_data = 12'h000;
			{8'd54, 8'd81}: color_data = 12'h000;
			{8'd54, 8'd85}: color_data = 12'h000;
			{8'd54, 8'd86}: color_data = 12'h112;
			{8'd54, 8'd87}: color_data = 12'h479;
			{8'd54, 8'd88}: color_data = 12'h49b;
			{8'd54, 8'd89}: color_data = 12'h48a;
			{8'd54, 8'd90}: color_data = 12'h48a;
			{8'd54, 8'd91}: color_data = 12'h48a;
			{8'd54, 8'd92}: color_data = 12'h48a;
			{8'd54, 8'd93}: color_data = 12'h48a;
			{8'd54, 8'd94}: color_data = 12'h48a;
			{8'd54, 8'd95}: color_data = 12'h48a;
			{8'd54, 8'd96}: color_data = 12'h48a;
			{8'd54, 8'd97}: color_data = 12'h48a;
			{8'd54, 8'd98}: color_data = 12'h48a;
			{8'd54, 8'd99}: color_data = 12'h48a;
			{8'd54, 8'd100}: color_data = 12'h48a;
			{8'd54, 8'd101}: color_data = 12'h48a;
			{8'd54, 8'd102}: color_data = 12'h48a;
			{8'd54, 8'd103}: color_data = 12'h48a;
			{8'd54, 8'd104}: color_data = 12'h48a;
			{8'd54, 8'd105}: color_data = 12'h48a;
			{8'd54, 8'd106}: color_data = 12'h48a;
			{8'd54, 8'd107}: color_data = 12'h48a;
			{8'd54, 8'd108}: color_data = 12'h48a;
			{8'd54, 8'd109}: color_data = 12'h49b;
			{8'd54, 8'd110}: color_data = 12'h367;
			{8'd54, 8'd111}: color_data = 12'h632;
			{8'd54, 8'd112}: color_data = 12'h942;
			{8'd54, 8'd113}: color_data = 12'h732;
			{8'd54, 8'd114}: color_data = 12'h742;
			{8'd54, 8'd115}: color_data = 12'hd95;
			{8'd54, 8'd116}: color_data = 12'hfb6;
			{8'd54, 8'd117}: color_data = 12'hfb6;
			{8'd54, 8'd118}: color_data = 12'hfb6;
			{8'd54, 8'd119}: color_data = 12'hfb6;
			{8'd54, 8'd120}: color_data = 12'hfb6;
			{8'd54, 8'd121}: color_data = 12'hfb6;
			{8'd54, 8'd122}: color_data = 12'hfb6;
			{8'd54, 8'd123}: color_data = 12'hfb6;
			{8'd54, 8'd124}: color_data = 12'hfb6;
			{8'd54, 8'd125}: color_data = 12'hfb6;
			{8'd54, 8'd126}: color_data = 12'hfb6;
			{8'd54, 8'd127}: color_data = 12'hfb6;
			{8'd54, 8'd128}: color_data = 12'hfa6;
			{8'd54, 8'd129}: color_data = 12'ha74;
			{8'd54, 8'd130}: color_data = 12'ha74;
			{8'd54, 8'd131}: color_data = 12'hea6;
			{8'd54, 8'd132}: color_data = 12'hfb6;
			{8'd54, 8'd133}: color_data = 12'hfb6;
			{8'd54, 8'd134}: color_data = 12'ha74;
			{8'd54, 8'd135}: color_data = 12'h211;
			{8'd55, 8'd28}: color_data = 12'hfc6;
			{8'd55, 8'd29}: color_data = 12'hfc4;
			{8'd55, 8'd30}: color_data = 12'hfc5;
			{8'd55, 8'd86}: color_data = 12'h000;
			{8'd55, 8'd87}: color_data = 12'h123;
			{8'd55, 8'd88}: color_data = 12'h479;
			{8'd55, 8'd89}: color_data = 12'h49b;
			{8'd55, 8'd90}: color_data = 12'h48a;
			{8'd55, 8'd91}: color_data = 12'h48a;
			{8'd55, 8'd92}: color_data = 12'h48a;
			{8'd55, 8'd93}: color_data = 12'h48a;
			{8'd55, 8'd94}: color_data = 12'h48a;
			{8'd55, 8'd95}: color_data = 12'h48a;
			{8'd55, 8'd96}: color_data = 12'h48a;
			{8'd55, 8'd97}: color_data = 12'h48a;
			{8'd55, 8'd98}: color_data = 12'h48a;
			{8'd55, 8'd99}: color_data = 12'h48a;
			{8'd55, 8'd100}: color_data = 12'h48a;
			{8'd55, 8'd101}: color_data = 12'h48a;
			{8'd55, 8'd102}: color_data = 12'h48a;
			{8'd55, 8'd103}: color_data = 12'h48a;
			{8'd55, 8'd104}: color_data = 12'h48a;
			{8'd55, 8'd105}: color_data = 12'h48a;
			{8'd55, 8'd106}: color_data = 12'h48a;
			{8'd55, 8'd107}: color_data = 12'h48a;
			{8'd55, 8'd108}: color_data = 12'h48a;
			{8'd55, 8'd109}: color_data = 12'h48a;
			{8'd55, 8'd110}: color_data = 12'h49b;
			{8'd55, 8'd111}: color_data = 12'h367;
			{8'd55, 8'd112}: color_data = 12'h532;
			{8'd55, 8'd113}: color_data = 12'h842;
			{8'd55, 8'd114}: color_data = 12'h842;
			{8'd55, 8'd115}: color_data = 12'h632;
			{8'd55, 8'd116}: color_data = 12'ha74;
			{8'd55, 8'd117}: color_data = 12'hfb6;
			{8'd55, 8'd118}: color_data = 12'hfb6;
			{8'd55, 8'd119}: color_data = 12'hfb6;
			{8'd55, 8'd120}: color_data = 12'hfb6;
			{8'd55, 8'd121}: color_data = 12'hfb6;
			{8'd55, 8'd122}: color_data = 12'hfb6;
			{8'd55, 8'd123}: color_data = 12'hfb6;
			{8'd55, 8'd124}: color_data = 12'hfb6;
			{8'd55, 8'd125}: color_data = 12'hfb6;
			{8'd55, 8'd126}: color_data = 12'hfb6;
			{8'd55, 8'd127}: color_data = 12'hfb6;
			{8'd55, 8'd128}: color_data = 12'hd95;
			{8'd55, 8'd129}: color_data = 12'ha74;
			{8'd55, 8'd130}: color_data = 12'ha74;
			{8'd55, 8'd131}: color_data = 12'hfb6;
			{8'd55, 8'd132}: color_data = 12'hfb6;
			{8'd55, 8'd133}: color_data = 12'hfb6;
			{8'd55, 8'd134}: color_data = 12'hfb7;
			{8'd55, 8'd135}: color_data = 12'hb84;
			{8'd55, 8'd136}: color_data = 12'h100;
			{8'd56, 8'd87}: color_data = 12'h000;
			{8'd56, 8'd88}: color_data = 12'h123;
			{8'd56, 8'd89}: color_data = 12'h379;
			{8'd56, 8'd90}: color_data = 12'h49b;
			{8'd56, 8'd91}: color_data = 12'h48a;
			{8'd56, 8'd92}: color_data = 12'h48a;
			{8'd56, 8'd93}: color_data = 12'h48a;
			{8'd56, 8'd94}: color_data = 12'h48a;
			{8'd56, 8'd95}: color_data = 12'h48a;
			{8'd56, 8'd96}: color_data = 12'h48a;
			{8'd56, 8'd97}: color_data = 12'h48a;
			{8'd56, 8'd98}: color_data = 12'h48a;
			{8'd56, 8'd99}: color_data = 12'h48a;
			{8'd56, 8'd100}: color_data = 12'h48a;
			{8'd56, 8'd101}: color_data = 12'h48a;
			{8'd56, 8'd102}: color_data = 12'h48a;
			{8'd56, 8'd103}: color_data = 12'h48a;
			{8'd56, 8'd104}: color_data = 12'h48a;
			{8'd56, 8'd105}: color_data = 12'h48a;
			{8'd56, 8'd106}: color_data = 12'h48a;
			{8'd56, 8'd107}: color_data = 12'h48a;
			{8'd56, 8'd108}: color_data = 12'h48a;
			{8'd56, 8'd109}: color_data = 12'h48b;
			{8'd56, 8'd110}: color_data = 12'h49b;
			{8'd56, 8'd111}: color_data = 12'h59b;
			{8'd56, 8'd112}: color_data = 12'h379;
			{8'd56, 8'd113}: color_data = 12'h443;
			{8'd56, 8'd114}: color_data = 12'h742;
			{8'd56, 8'd115}: color_data = 12'h842;
			{8'd56, 8'd116}: color_data = 12'h732;
			{8'd56, 8'd117}: color_data = 12'h642;
			{8'd56, 8'd118}: color_data = 12'hc85;
			{8'd56, 8'd119}: color_data = 12'hfb6;
			{8'd56, 8'd120}: color_data = 12'hfb6;
			{8'd56, 8'd121}: color_data = 12'hfb6;
			{8'd56, 8'd122}: color_data = 12'hfb6;
			{8'd56, 8'd123}: color_data = 12'hfb6;
			{8'd56, 8'd124}: color_data = 12'hfb6;
			{8'd56, 8'd125}: color_data = 12'hfb6;
			{8'd56, 8'd126}: color_data = 12'hfb6;
			{8'd56, 8'd127}: color_data = 12'hfb6;
			{8'd56, 8'd128}: color_data = 12'ha74;
			{8'd56, 8'd129}: color_data = 12'ha74;
			{8'd56, 8'd130}: color_data = 12'hc85;
			{8'd56, 8'd131}: color_data = 12'hfb6;
			{8'd56, 8'd132}: color_data = 12'hfb6;
			{8'd56, 8'd133}: color_data = 12'hfb6;
			{8'd56, 8'd134}: color_data = 12'hfb6;
			{8'd56, 8'd135}: color_data = 12'hfb7;
			{8'd56, 8'd136}: color_data = 12'h863;
			{8'd56, 8'd137}: color_data = 12'h000;
			{8'd57, 8'd13}: color_data = 12'hfc4;
			{8'd57, 8'd14}: color_data = 12'hfc4;
			{8'd57, 8'd15}: color_data = 12'heb2;
			{8'd57, 8'd16}: color_data = 12'heb4;
			{8'd57, 8'd17}: color_data = 12'hfc6;
			{8'd57, 8'd89}: color_data = 12'h112;
			{8'd57, 8'd90}: color_data = 12'h367;
			{8'd57, 8'd91}: color_data = 12'h49b;
			{8'd57, 8'd92}: color_data = 12'h48b;
			{8'd57, 8'd93}: color_data = 12'h48a;
			{8'd57, 8'd94}: color_data = 12'h48a;
			{8'd57, 8'd95}: color_data = 12'h48a;
			{8'd57, 8'd96}: color_data = 12'h48a;
			{8'd57, 8'd97}: color_data = 12'h48a;
			{8'd57, 8'd98}: color_data = 12'h48a;
			{8'd57, 8'd99}: color_data = 12'h48a;
			{8'd57, 8'd100}: color_data = 12'h48a;
			{8'd57, 8'd101}: color_data = 12'h48a;
			{8'd57, 8'd102}: color_data = 12'h48a;
			{8'd57, 8'd103}: color_data = 12'h48a;
			{8'd57, 8'd104}: color_data = 12'h48a;
			{8'd57, 8'd105}: color_data = 12'h48a;
			{8'd57, 8'd106}: color_data = 12'h48a;
			{8'd57, 8'd107}: color_data = 12'h48b;
			{8'd57, 8'd108}: color_data = 12'h48b;
			{8'd57, 8'd109}: color_data = 12'h479;
			{8'd57, 8'd110}: color_data = 12'h368;
			{8'd57, 8'd111}: color_data = 12'h257;
			{8'd57, 8'd112}: color_data = 12'h257;
			{8'd57, 8'd113}: color_data = 12'h146;
			{8'd57, 8'd114}: color_data = 12'h023;
			{8'd57, 8'd115}: color_data = 12'h322;
			{8'd57, 8'd116}: color_data = 12'h842;
			{8'd57, 8'd117}: color_data = 12'h842;
			{8'd57, 8'd118}: color_data = 12'h632;
			{8'd57, 8'd119}: color_data = 12'h753;
			{8'd57, 8'd120}: color_data = 12'hc85;
			{8'd57, 8'd121}: color_data = 12'hfb6;
			{8'd57, 8'd122}: color_data = 12'hfb6;
			{8'd57, 8'd123}: color_data = 12'hfb6;
			{8'd57, 8'd124}: color_data = 12'hfb6;
			{8'd57, 8'd125}: color_data = 12'hfb6;
			{8'd57, 8'd126}: color_data = 12'hfb6;
			{8'd57, 8'd127}: color_data = 12'hd95;
			{8'd57, 8'd128}: color_data = 12'h964;
			{8'd57, 8'd129}: color_data = 12'h974;
			{8'd57, 8'd130}: color_data = 12'hfb6;
			{8'd57, 8'd131}: color_data = 12'hfb6;
			{8'd57, 8'd132}: color_data = 12'hfb6;
			{8'd57, 8'd133}: color_data = 12'hfb6;
			{8'd57, 8'd134}: color_data = 12'hfb6;
			{8'd57, 8'd135}: color_data = 12'hfb6;
			{8'd57, 8'd136}: color_data = 12'hd95;
			{8'd57, 8'd137}: color_data = 12'h211;
			{8'd58, 8'd12}: color_data = 12'hfd5;
			{8'd58, 8'd13}: color_data = 12'hfc5;
			{8'd58, 8'd14}: color_data = 12'hfc5;
			{8'd58, 8'd15}: color_data = 12'hfc5;
			{8'd58, 8'd16}: color_data = 12'hfc4;
			{8'd58, 8'd17}: color_data = 12'hfc5;
			{8'd58, 8'd18}: color_data = 12'hfc5;
			{8'd58, 8'd19}: color_data = 12'hec5;
			{8'd58, 8'd90}: color_data = 12'h000;
			{8'd58, 8'd91}: color_data = 12'h246;
			{8'd58, 8'd92}: color_data = 12'h48a;
			{8'd58, 8'd93}: color_data = 12'h49b;
			{8'd58, 8'd94}: color_data = 12'h48b;
			{8'd58, 8'd95}: color_data = 12'h48a;
			{8'd58, 8'd96}: color_data = 12'h48a;
			{8'd58, 8'd97}: color_data = 12'h48a;
			{8'd58, 8'd98}: color_data = 12'h48a;
			{8'd58, 8'd99}: color_data = 12'h48a;
			{8'd58, 8'd100}: color_data = 12'h48a;
			{8'd58, 8'd101}: color_data = 12'h48a;
			{8'd58, 8'd102}: color_data = 12'h48a;
			{8'd58, 8'd103}: color_data = 12'h48a;
			{8'd58, 8'd104}: color_data = 12'h48a;
			{8'd58, 8'd105}: color_data = 12'h48a;
			{8'd58, 8'd106}: color_data = 12'h48b;
			{8'd58, 8'd107}: color_data = 12'h479;
			{8'd58, 8'd108}: color_data = 12'h146;
			{8'd58, 8'd109}: color_data = 12'h047;
			{8'd58, 8'd110}: color_data = 12'h059;
			{8'd58, 8'd111}: color_data = 12'h05a;
			{8'd58, 8'd112}: color_data = 12'h05a;
			{8'd58, 8'd113}: color_data = 12'h05a;
			{8'd58, 8'd114}: color_data = 12'h037;
			{8'd58, 8'd115}: color_data = 12'h059;
			{8'd58, 8'd116}: color_data = 12'h333;
			{8'd58, 8'd117}: color_data = 12'h842;
			{8'd58, 8'd118}: color_data = 12'h942;
			{8'd58, 8'd119}: color_data = 12'h842;
			{8'd58, 8'd120}: color_data = 12'h632;
			{8'd58, 8'd121}: color_data = 12'h742;
			{8'd58, 8'd122}: color_data = 12'h963;
			{8'd58, 8'd123}: color_data = 12'hc85;
			{8'd58, 8'd124}: color_data = 12'hea6;
			{8'd58, 8'd125}: color_data = 12'hfb6;
			{8'd58, 8'd126}: color_data = 12'hfa6;
			{8'd58, 8'd127}: color_data = 12'h964;
			{8'd58, 8'd128}: color_data = 12'h964;
			{8'd58, 8'd129}: color_data = 12'hd95;
			{8'd58, 8'd130}: color_data = 12'hfb6;
			{8'd58, 8'd131}: color_data = 12'hfb6;
			{8'd58, 8'd132}: color_data = 12'hfb6;
			{8'd58, 8'd133}: color_data = 12'hfb6;
			{8'd58, 8'd134}: color_data = 12'hfb6;
			{8'd58, 8'd135}: color_data = 12'hfb6;
			{8'd58, 8'd136}: color_data = 12'hfb6;
			{8'd58, 8'd137}: color_data = 12'h653;
			{8'd59, 8'd12}: color_data = 12'hfc5;
			{8'd59, 8'd13}: color_data = 12'hfc5;
			{8'd59, 8'd14}: color_data = 12'hfc4;
			{8'd59, 8'd15}: color_data = 12'hfb2;
			{8'd59, 8'd16}: color_data = 12'hfc4;
			{8'd59, 8'd17}: color_data = 12'hfc5;
			{8'd59, 8'd18}: color_data = 12'hfc5;
			{8'd59, 8'd19}: color_data = 12'hfc4;
			{8'd59, 8'd20}: color_data = 12'hfc5;
			{8'd59, 8'd21}: color_data = 12'hfd5;
			{8'd59, 8'd91}: color_data = 12'h000;
			{8'd59, 8'd92}: color_data = 12'h123;
			{8'd59, 8'd93}: color_data = 12'h357;
			{8'd59, 8'd94}: color_data = 12'h48a;
			{8'd59, 8'd95}: color_data = 12'h48b;
			{8'd59, 8'd96}: color_data = 12'h49b;
			{8'd59, 8'd97}: color_data = 12'h48b;
			{8'd59, 8'd98}: color_data = 12'h48a;
			{8'd59, 8'd99}: color_data = 12'h48a;
			{8'd59, 8'd100}: color_data = 12'h48a;
			{8'd59, 8'd101}: color_data = 12'h48a;
			{8'd59, 8'd102}: color_data = 12'h48a;
			{8'd59, 8'd103}: color_data = 12'h48a;
			{8'd59, 8'd104}: color_data = 12'h48a;
			{8'd59, 8'd105}: color_data = 12'h48b;
			{8'd59, 8'd106}: color_data = 12'h368;
			{8'd59, 8'd107}: color_data = 12'h047;
			{8'd59, 8'd108}: color_data = 12'h05a;
			{8'd59, 8'd109}: color_data = 12'h06b;
			{8'd59, 8'd110}: color_data = 12'h06b;
			{8'd59, 8'd111}: color_data = 12'h06b;
			{8'd59, 8'd112}: color_data = 12'h06b;
			{8'd59, 8'd113}: color_data = 12'h06b;
			{8'd59, 8'd114}: color_data = 12'h059;
			{8'd59, 8'd115}: color_data = 12'h047;
			{8'd59, 8'd116}: color_data = 12'h06a;
			{8'd59, 8'd117}: color_data = 12'h146;
			{8'd59, 8'd118}: color_data = 12'h432;
			{8'd59, 8'd119}: color_data = 12'h842;
			{8'd59, 8'd120}: color_data = 12'h942;
			{8'd59, 8'd121}: color_data = 12'h842;
			{8'd59, 8'd122}: color_data = 12'h742;
			{8'd59, 8'd123}: color_data = 12'h632;
			{8'd59, 8'd124}: color_data = 12'h632;
			{8'd59, 8'd125}: color_data = 12'h742;
			{8'd59, 8'd126}: color_data = 12'h532;
			{8'd59, 8'd127}: color_data = 12'h753;
			{8'd59, 8'd128}: color_data = 12'h863;
			{8'd59, 8'd129}: color_data = 12'hfb6;
			{8'd59, 8'd130}: color_data = 12'hfb6;
			{8'd59, 8'd131}: color_data = 12'hfb6;
			{8'd59, 8'd132}: color_data = 12'hfb6;
			{8'd59, 8'd133}: color_data = 12'hfb6;
			{8'd59, 8'd134}: color_data = 12'hfb6;
			{8'd59, 8'd135}: color_data = 12'hfb6;
			{8'd59, 8'd136}: color_data = 12'hfb7;
			{8'd59, 8'd137}: color_data = 12'h963;
			{8'd59, 8'd138}: color_data = 12'h000;
			{8'd60, 8'd12}: color_data = 12'hfc4;
			{8'd60, 8'd13}: color_data = 12'hfc5;
			{8'd60, 8'd14}: color_data = 12'heb2;
			{8'd60, 8'd15}: color_data = 12'hd90;
			{8'd60, 8'd16}: color_data = 12'hd90;
			{8'd60, 8'd17}: color_data = 12'hea2;
			{8'd60, 8'd18}: color_data = 12'hfc4;
			{8'd60, 8'd19}: color_data = 12'hfc5;
			{8'd60, 8'd20}: color_data = 12'hfc5;
			{8'd60, 8'd21}: color_data = 12'hfc5;
			{8'd60, 8'd22}: color_data = 12'hfc5;
			{8'd60, 8'd23}: color_data = 12'hfc7;
			{8'd60, 8'd93}: color_data = 12'h000;
			{8'd60, 8'd94}: color_data = 12'h122;
			{8'd60, 8'd95}: color_data = 12'h134;
			{8'd60, 8'd96}: color_data = 12'h235;
			{8'd60, 8'd97}: color_data = 12'h378;
			{8'd60, 8'd98}: color_data = 12'h49b;
			{8'd60, 8'd99}: color_data = 12'h48a;
			{8'd60, 8'd100}: color_data = 12'h48a;
			{8'd60, 8'd101}: color_data = 12'h48a;
			{8'd60, 8'd102}: color_data = 12'h48a;
			{8'd60, 8'd103}: color_data = 12'h48a;
			{8'd60, 8'd104}: color_data = 12'h48b;
			{8'd60, 8'd105}: color_data = 12'h479;
			{8'd60, 8'd106}: color_data = 12'h047;
			{8'd60, 8'd107}: color_data = 12'h06b;
			{8'd60, 8'd108}: color_data = 12'h06b;
			{8'd60, 8'd109}: color_data = 12'h06b;
			{8'd60, 8'd110}: color_data = 12'h06b;
			{8'd60, 8'd111}: color_data = 12'h06b;
			{8'd60, 8'd112}: color_data = 12'h06b;
			{8'd60, 8'd113}: color_data = 12'h06b;
			{8'd60, 8'd114}: color_data = 12'h06b;
			{8'd60, 8'd115}: color_data = 12'h048;
			{8'd60, 8'd116}: color_data = 12'h047;
			{8'd60, 8'd117}: color_data = 12'h06b;
			{8'd60, 8'd118}: color_data = 12'h05a;
			{8'd60, 8'd119}: color_data = 12'h146;
			{8'd60, 8'd120}: color_data = 12'h432;
			{8'd60, 8'd121}: color_data = 12'h732;
			{8'd60, 8'd122}: color_data = 12'h842;
			{8'd60, 8'd123}: color_data = 12'h843;
			{8'd60, 8'd124}: color_data = 12'h842;
			{8'd60, 8'd125}: color_data = 12'h842;
			{8'd60, 8'd126}: color_data = 12'h632;
			{8'd60, 8'd127}: color_data = 12'h964;
			{8'd60, 8'd128}: color_data = 12'hd95;
			{8'd60, 8'd129}: color_data = 12'ha74;
			{8'd60, 8'd130}: color_data = 12'hfb6;
			{8'd60, 8'd131}: color_data = 12'hfb6;
			{8'd60, 8'd132}: color_data = 12'hfb6;
			{8'd60, 8'd133}: color_data = 12'hfb6;
			{8'd60, 8'd134}: color_data = 12'hfb6;
			{8'd60, 8'd135}: color_data = 12'hfb6;
			{8'd60, 8'd136}: color_data = 12'hfb7;
			{8'd60, 8'd137}: color_data = 12'h964;
			{8'd60, 8'd138}: color_data = 12'h000;
			{8'd61, 8'd11}: color_data = 12'hfc5;
			{8'd61, 8'd12}: color_data = 12'hfc5;
			{8'd61, 8'd13}: color_data = 12'hfc5;
			{8'd61, 8'd14}: color_data = 12'hea1;
			{8'd61, 8'd15}: color_data = 12'hd90;
			{8'd61, 8'd16}: color_data = 12'hd90;
			{8'd61, 8'd17}: color_data = 12'hd90;
			{8'd61, 8'd18}: color_data = 12'hd90;
			{8'd61, 8'd19}: color_data = 12'hea1;
			{8'd61, 8'd20}: color_data = 12'hfc4;
			{8'd61, 8'd21}: color_data = 12'hfc5;
			{8'd61, 8'd22}: color_data = 12'hfc5;
			{8'd61, 8'd23}: color_data = 12'hfc4;
			{8'd61, 8'd24}: color_data = 12'hfc5;
			{8'd61, 8'd25}: color_data = 12'hfc5;
			{8'd61, 8'd97}: color_data = 12'h012;
			{8'd61, 8'd98}: color_data = 12'h368;
			{8'd61, 8'd99}: color_data = 12'h49b;
			{8'd61, 8'd100}: color_data = 12'h48b;
			{8'd61, 8'd101}: color_data = 12'h48a;
			{8'd61, 8'd102}: color_data = 12'h48a;
			{8'd61, 8'd103}: color_data = 12'h48a;
			{8'd61, 8'd104}: color_data = 12'h49b;
			{8'd61, 8'd105}: color_data = 12'h367;
			{8'd61, 8'd106}: color_data = 12'h059;
			{8'd61, 8'd107}: color_data = 12'h06b;
			{8'd61, 8'd108}: color_data = 12'h06b;
			{8'd61, 8'd109}: color_data = 12'h06b;
			{8'd61, 8'd110}: color_data = 12'h06b;
			{8'd61, 8'd111}: color_data = 12'h06b;
			{8'd61, 8'd112}: color_data = 12'h06b;
			{8'd61, 8'd113}: color_data = 12'h06b;
			{8'd61, 8'd114}: color_data = 12'h06b;
			{8'd61, 8'd115}: color_data = 12'h06b;
			{8'd61, 8'd116}: color_data = 12'h048;
			{8'd61, 8'd117}: color_data = 12'h047;
			{8'd61, 8'd118}: color_data = 12'h06b;
			{8'd61, 8'd119}: color_data = 12'h06b;
			{8'd61, 8'd120}: color_data = 12'h059;
			{8'd61, 8'd121}: color_data = 12'h222;
			{8'd61, 8'd122}: color_data = 12'h531;
			{8'd61, 8'd123}: color_data = 12'h842;
			{8'd61, 8'd124}: color_data = 12'h842;
			{8'd61, 8'd125}: color_data = 12'h842;
			{8'd61, 8'd126}: color_data = 12'h843;
			{8'd61, 8'd127}: color_data = 12'h632;
			{8'd61, 8'd128}: color_data = 12'ha74;
			{8'd61, 8'd129}: color_data = 12'hd95;
			{8'd61, 8'd130}: color_data = 12'h974;
			{8'd61, 8'd131}: color_data = 12'hd95;
			{8'd61, 8'd132}: color_data = 12'hfb6;
			{8'd61, 8'd133}: color_data = 12'hfb6;
			{8'd61, 8'd134}: color_data = 12'hfb6;
			{8'd61, 8'd135}: color_data = 12'hfb6;
			{8'd61, 8'd136}: color_data = 12'hfb6;
			{8'd61, 8'd137}: color_data = 12'h642;
			{8'd62, 8'd11}: color_data = 12'hfc5;
			{8'd62, 8'd12}: color_data = 12'hfc5;
			{8'd62, 8'd13}: color_data = 12'hfc4;
			{8'd62, 8'd14}: color_data = 12'hd90;
			{8'd62, 8'd15}: color_data = 12'hd90;
			{8'd62, 8'd16}: color_data = 12'hd90;
			{8'd62, 8'd17}: color_data = 12'hd90;
			{8'd62, 8'd18}: color_data = 12'hd90;
			{8'd62, 8'd19}: color_data = 12'hd90;
			{8'd62, 8'd20}: color_data = 12'hd90;
			{8'd62, 8'd21}: color_data = 12'hea1;
			{8'd62, 8'd22}: color_data = 12'hfc4;
			{8'd62, 8'd23}: color_data = 12'hfc5;
			{8'd62, 8'd24}: color_data = 12'hfc5;
			{8'd62, 8'd25}: color_data = 12'hfc5;
			{8'd62, 8'd26}: color_data = 12'hfc5;
			{8'd62, 8'd27}: color_data = 12'heb5;
			{8'd62, 8'd98}: color_data = 12'h001;
			{8'd62, 8'd99}: color_data = 12'h256;
			{8'd62, 8'd100}: color_data = 12'h48a;
			{8'd62, 8'd101}: color_data = 12'h49b;
			{8'd62, 8'd102}: color_data = 12'h48b;
			{8'd62, 8'd103}: color_data = 12'h48a;
			{8'd62, 8'd104}: color_data = 12'h49b;
			{8'd62, 8'd105}: color_data = 12'h257;
			{8'd62, 8'd106}: color_data = 12'h05a;
			{8'd62, 8'd107}: color_data = 12'h06b;
			{8'd62, 8'd108}: color_data = 12'h06b;
			{8'd62, 8'd109}: color_data = 12'h06b;
			{8'd62, 8'd110}: color_data = 12'h06b;
			{8'd62, 8'd111}: color_data = 12'h06b;
			{8'd62, 8'd112}: color_data = 12'h06b;
			{8'd62, 8'd113}: color_data = 12'h06b;
			{8'd62, 8'd114}: color_data = 12'h06b;
			{8'd62, 8'd115}: color_data = 12'h06b;
			{8'd62, 8'd116}: color_data = 12'h06b;
			{8'd62, 8'd117}: color_data = 12'h06a;
			{8'd62, 8'd118}: color_data = 12'h06b;
			{8'd62, 8'd119}: color_data = 12'h06b;
			{8'd62, 8'd120}: color_data = 12'h06b;
			{8'd62, 8'd121}: color_data = 12'h059;
			{8'd62, 8'd122}: color_data = 12'h432;
			{8'd62, 8'd123}: color_data = 12'h842;
			{8'd62, 8'd124}: color_data = 12'h843;
			{8'd62, 8'd125}: color_data = 12'h842;
			{8'd62, 8'd126}: color_data = 12'h842;
			{8'd62, 8'd127}: color_data = 12'h842;
			{8'd62, 8'd128}: color_data = 12'h632;
			{8'd62, 8'd129}: color_data = 12'h853;
			{8'd62, 8'd130}: color_data = 12'hb84;
			{8'd62, 8'd131}: color_data = 12'h974;
			{8'd62, 8'd132}: color_data = 12'ha74;
			{8'd62, 8'd133}: color_data = 12'hd95;
			{8'd62, 8'd134}: color_data = 12'hea6;
			{8'd62, 8'd135}: color_data = 12'hda5;
			{8'd62, 8'd136}: color_data = 12'ha74;
			{8'd62, 8'd137}: color_data = 12'h110;
			{8'd63, 8'd11}: color_data = 12'hfc5;
			{8'd63, 8'd12}: color_data = 12'hfc5;
			{8'd63, 8'd13}: color_data = 12'hfc4;
			{8'd63, 8'd14}: color_data = 12'hea1;
			{8'd63, 8'd15}: color_data = 12'hd90;
			{8'd63, 8'd16}: color_data = 12'hd90;
			{8'd63, 8'd17}: color_data = 12'hd90;
			{8'd63, 8'd18}: color_data = 12'hd90;
			{8'd63, 8'd19}: color_data = 12'hd90;
			{8'd63, 8'd20}: color_data = 12'hd90;
			{8'd63, 8'd21}: color_data = 12'hd90;
			{8'd63, 8'd22}: color_data = 12'hd90;
			{8'd63, 8'd23}: color_data = 12'hea1;
			{8'd63, 8'd24}: color_data = 12'hfc4;
			{8'd63, 8'd25}: color_data = 12'hfc5;
			{8'd63, 8'd26}: color_data = 12'hfc5;
			{8'd63, 8'd27}: color_data = 12'hfc5;
			{8'd63, 8'd28}: color_data = 12'hfc5;
			{8'd63, 8'd92}: color_data = 12'h000;
			{8'd63, 8'd93}: color_data = 12'h100;
			{8'd63, 8'd94}: color_data = 12'h400;
			{8'd63, 8'd95}: color_data = 12'h601;
			{8'd63, 8'd96}: color_data = 12'h500;
			{8'd63, 8'd97}: color_data = 12'h300;
			{8'd63, 8'd98}: color_data = 12'h000;
			{8'd63, 8'd99}: color_data = 12'h000;
			{8'd63, 8'd100}: color_data = 12'h134;
			{8'd63, 8'd101}: color_data = 12'h368;
			{8'd63, 8'd102}: color_data = 12'h48a;
			{8'd63, 8'd103}: color_data = 12'h49b;
			{8'd63, 8'd104}: color_data = 12'h59b;
			{8'd63, 8'd105}: color_data = 12'h368;
			{8'd63, 8'd106}: color_data = 12'h059;
			{8'd63, 8'd107}: color_data = 12'h06b;
			{8'd63, 8'd108}: color_data = 12'h06b;
			{8'd63, 8'd109}: color_data = 12'h06b;
			{8'd63, 8'd110}: color_data = 12'h06b;
			{8'd63, 8'd111}: color_data = 12'h06b;
			{8'd63, 8'd112}: color_data = 12'h06b;
			{8'd63, 8'd113}: color_data = 12'h06b;
			{8'd63, 8'd114}: color_data = 12'h06b;
			{8'd63, 8'd115}: color_data = 12'h06b;
			{8'd63, 8'd116}: color_data = 12'h06b;
			{8'd63, 8'd117}: color_data = 12'h06b;
			{8'd63, 8'd118}: color_data = 12'h06b;
			{8'd63, 8'd119}: color_data = 12'h06b;
			{8'd63, 8'd120}: color_data = 12'h06b;
			{8'd63, 8'd121}: color_data = 12'h06b;
			{8'd63, 8'd122}: color_data = 12'h059;
			{8'd63, 8'd123}: color_data = 12'h432;
			{8'd63, 8'd124}: color_data = 12'h842;
			{8'd63, 8'd125}: color_data = 12'h843;
			{8'd63, 8'd126}: color_data = 12'h842;
			{8'd63, 8'd127}: color_data = 12'h842;
			{8'd63, 8'd128}: color_data = 12'h843;
			{8'd63, 8'd129}: color_data = 12'h842;
			{8'd63, 8'd130}: color_data = 12'h632;
			{8'd63, 8'd131}: color_data = 12'h742;
			{8'd63, 8'd132}: color_data = 12'h742;
			{8'd63, 8'd133}: color_data = 12'h642;
			{8'd63, 8'd134}: color_data = 12'h753;
			{8'd63, 8'd135}: color_data = 12'h863;
			{8'd63, 8'd136}: color_data = 12'h210;
			{8'd64, 8'd11}: color_data = 12'hfc4;
			{8'd64, 8'd12}: color_data = 12'hfc4;
			{8'd64, 8'd13}: color_data = 12'hfc5;
			{8'd64, 8'd14}: color_data = 12'hfc5;
			{8'd64, 8'd15}: color_data = 12'hfb4;
			{8'd64, 8'd16}: color_data = 12'hea1;
			{8'd64, 8'd17}: color_data = 12'hd90;
			{8'd64, 8'd18}: color_data = 12'hd90;
			{8'd64, 8'd19}: color_data = 12'hd90;
			{8'd64, 8'd20}: color_data = 12'hd90;
			{8'd64, 8'd21}: color_data = 12'hd90;
			{8'd64, 8'd22}: color_data = 12'hd90;
			{8'd64, 8'd23}: color_data = 12'hd90;
			{8'd64, 8'd24}: color_data = 12'hd90;
			{8'd64, 8'd25}: color_data = 12'hea1;
			{8'd64, 8'd26}: color_data = 12'hfb4;
			{8'd64, 8'd27}: color_data = 12'hfc5;
			{8'd64, 8'd28}: color_data = 12'hfc5;
			{8'd64, 8'd29}: color_data = 12'hfc5;
			{8'd64, 8'd91}: color_data = 12'h000;
			{8'd64, 8'd92}: color_data = 12'h601;
			{8'd64, 8'd93}: color_data = 12'hb11;
			{8'd64, 8'd94}: color_data = 12'he12;
			{8'd64, 8'd95}: color_data = 12'hf12;
			{8'd64, 8'd96}: color_data = 12'hf12;
			{8'd64, 8'd97}: color_data = 12'hd12;
			{8'd64, 8'd98}: color_data = 12'h911;
			{8'd64, 8'd99}: color_data = 12'h200;
			{8'd64, 8'd101}: color_data = 12'h000;
			{8'd64, 8'd102}: color_data = 12'h134;
			{8'd64, 8'd103}: color_data = 12'h246;
			{8'd64, 8'd104}: color_data = 12'h357;
			{8'd64, 8'd105}: color_data = 12'h246;
			{8'd64, 8'd106}: color_data = 12'h047;
			{8'd64, 8'd107}: color_data = 12'h06b;
			{8'd64, 8'd108}: color_data = 12'h06b;
			{8'd64, 8'd109}: color_data = 12'h06b;
			{8'd64, 8'd110}: color_data = 12'h06b;
			{8'd64, 8'd111}: color_data = 12'h06b;
			{8'd64, 8'd112}: color_data = 12'h06b;
			{8'd64, 8'd113}: color_data = 12'h06b;
			{8'd64, 8'd114}: color_data = 12'h06b;
			{8'd64, 8'd115}: color_data = 12'h06b;
			{8'd64, 8'd116}: color_data = 12'h06b;
			{8'd64, 8'd117}: color_data = 12'h06b;
			{8'd64, 8'd118}: color_data = 12'h06b;
			{8'd64, 8'd119}: color_data = 12'h06b;
			{8'd64, 8'd120}: color_data = 12'h06b;
			{8'd64, 8'd121}: color_data = 12'h06b;
			{8'd64, 8'd122}: color_data = 12'h06b;
			{8'd64, 8'd123}: color_data = 12'h059;
			{8'd64, 8'd124}: color_data = 12'h234;
			{8'd64, 8'd125}: color_data = 12'h742;
			{8'd64, 8'd126}: color_data = 12'h842;
			{8'd64, 8'd127}: color_data = 12'h843;
			{8'd64, 8'd128}: color_data = 12'h842;
			{8'd64, 8'd129}: color_data = 12'h842;
			{8'd64, 8'd130}: color_data = 12'h843;
			{8'd64, 8'd131}: color_data = 12'h842;
			{8'd64, 8'd132}: color_data = 12'h842;
			{8'd64, 8'd133}: color_data = 12'h842;
			{8'd64, 8'd134}: color_data = 12'h632;
			{8'd64, 8'd135}: color_data = 12'h210;
			{8'd64, 8'd136}: color_data = 12'h000;
			{8'd65, 8'd12}: color_data = 12'hfc4;
			{8'd65, 8'd13}: color_data = 12'hfc5;
			{8'd65, 8'd14}: color_data = 12'hfc4;
			{8'd65, 8'd15}: color_data = 12'hfc5;
			{8'd65, 8'd16}: color_data = 12'hfc5;
			{8'd65, 8'd17}: color_data = 12'hfb4;
			{8'd65, 8'd18}: color_data = 12'hea1;
			{8'd65, 8'd19}: color_data = 12'hd90;
			{8'd65, 8'd20}: color_data = 12'hd90;
			{8'd65, 8'd21}: color_data = 12'hd90;
			{8'd65, 8'd22}: color_data = 12'hd90;
			{8'd65, 8'd23}: color_data = 12'hd90;
			{8'd65, 8'd24}: color_data = 12'hd90;
			{8'd65, 8'd25}: color_data = 12'hd90;
			{8'd65, 8'd26}: color_data = 12'hd90;
			{8'd65, 8'd27}: color_data = 12'hfb3;
			{8'd65, 8'd28}: color_data = 12'hfc5;
			{8'd65, 8'd29}: color_data = 12'hfc5;
			{8'd65, 8'd90}: color_data = 12'h000;
			{8'd65, 8'd91}: color_data = 12'h811;
			{8'd65, 8'd92}: color_data = 12'hf12;
			{8'd65, 8'd93}: color_data = 12'hf12;
			{8'd65, 8'd94}: color_data = 12'hf12;
			{8'd65, 8'd95}: color_data = 12'he12;
			{8'd65, 8'd96}: color_data = 12'he12;
			{8'd65, 8'd97}: color_data = 12'hf12;
			{8'd65, 8'd98}: color_data = 12'hf12;
			{8'd65, 8'd99}: color_data = 12'ha11;
			{8'd65, 8'd100}: color_data = 12'h000;
			{8'd65, 8'd103}: color_data = 12'h000;
			{8'd65, 8'd104}: color_data = 12'h000;
			{8'd65, 8'd105}: color_data = 12'h000;
			{8'd65, 8'd106}: color_data = 12'h035;
			{8'd65, 8'd107}: color_data = 12'h06b;
			{8'd65, 8'd108}: color_data = 12'h06b;
			{8'd65, 8'd109}: color_data = 12'h06b;
			{8'd65, 8'd110}: color_data = 12'h06b;
			{8'd65, 8'd111}: color_data = 12'h06b;
			{8'd65, 8'd112}: color_data = 12'h06b;
			{8'd65, 8'd113}: color_data = 12'h06b;
			{8'd65, 8'd114}: color_data = 12'h06b;
			{8'd65, 8'd115}: color_data = 12'h06b;
			{8'd65, 8'd116}: color_data = 12'h06b;
			{8'd65, 8'd117}: color_data = 12'h06b;
			{8'd65, 8'd118}: color_data = 12'h06b;
			{8'd65, 8'd119}: color_data = 12'h06b;
			{8'd65, 8'd120}: color_data = 12'h06b;
			{8'd65, 8'd121}: color_data = 12'h06b;
			{8'd65, 8'd122}: color_data = 12'h06b;
			{8'd65, 8'd123}: color_data = 12'h06b;
			{8'd65, 8'd124}: color_data = 12'h06b;
			{8'd65, 8'd125}: color_data = 12'h046;
			{8'd65, 8'd126}: color_data = 12'h433;
			{8'd65, 8'd127}: color_data = 12'h742;
			{8'd65, 8'd128}: color_data = 12'h842;
			{8'd65, 8'd129}: color_data = 12'h842;
			{8'd65, 8'd130}: color_data = 12'h843;
			{8'd65, 8'd131}: color_data = 12'h843;
			{8'd65, 8'd132}: color_data = 12'h843;
			{8'd65, 8'd133}: color_data = 12'h632;
			{8'd65, 8'd134}: color_data = 12'h210;
			{8'd65, 8'd135}: color_data = 12'h000;
			{8'd66, 8'd14}: color_data = 12'hec5;
			{8'd66, 8'd15}: color_data = 12'hfc6;
			{8'd66, 8'd16}: color_data = 12'hfc6;
			{8'd66, 8'd17}: color_data = 12'hfc5;
			{8'd66, 8'd18}: color_data = 12'hfc6;
			{8'd66, 8'd19}: color_data = 12'hea1;
			{8'd66, 8'd20}: color_data = 12'hd90;
			{8'd66, 8'd21}: color_data = 12'hd90;
			{8'd66, 8'd22}: color_data = 12'hd90;
			{8'd66, 8'd23}: color_data = 12'hd90;
			{8'd66, 8'd24}: color_data = 12'hd90;
			{8'd66, 8'd25}: color_data = 12'hd90;
			{8'd66, 8'd26}: color_data = 12'hd90;
			{8'd66, 8'd27}: color_data = 12'hfc4;
			{8'd66, 8'd28}: color_data = 12'hfc5;
			{8'd66, 8'd29}: color_data = 12'hfc5;
			{8'd66, 8'd57}: color_data = 12'h000;
			{8'd66, 8'd58}: color_data = 12'h200;
			{8'd66, 8'd59}: color_data = 12'h500;
			{8'd66, 8'd60}: color_data = 12'h400;
			{8'd66, 8'd61}: color_data = 12'h200;
			{8'd66, 8'd62}: color_data = 12'h000;
			{8'd66, 8'd89}: color_data = 12'h000;
			{8'd66, 8'd90}: color_data = 12'h801;
			{8'd66, 8'd91}: color_data = 12'hf12;
			{8'd66, 8'd92}: color_data = 12'hf11;
			{8'd66, 8'd93}: color_data = 12'he11;
			{8'd66, 8'd94}: color_data = 12'he11;
			{8'd66, 8'd95}: color_data = 12'he11;
			{8'd66, 8'd96}: color_data = 12'hf12;
			{8'd66, 8'd97}: color_data = 12'hf12;
			{8'd66, 8'd98}: color_data = 12'he12;
			{8'd66, 8'd99}: color_data = 12'he12;
			{8'd66, 8'd100}: color_data = 12'h500;
			{8'd66, 8'd106}: color_data = 12'h012;
			{8'd66, 8'd107}: color_data = 12'h059;
			{8'd66, 8'd108}: color_data = 12'h06b;
			{8'd66, 8'd109}: color_data = 12'h06b;
			{8'd66, 8'd110}: color_data = 12'h06b;
			{8'd66, 8'd111}: color_data = 12'h06b;
			{8'd66, 8'd112}: color_data = 12'h06b;
			{8'd66, 8'd113}: color_data = 12'h06b;
			{8'd66, 8'd114}: color_data = 12'h06b;
			{8'd66, 8'd115}: color_data = 12'h06b;
			{8'd66, 8'd116}: color_data = 12'h06b;
			{8'd66, 8'd117}: color_data = 12'h06b;
			{8'd66, 8'd118}: color_data = 12'h06b;
			{8'd66, 8'd119}: color_data = 12'h06b;
			{8'd66, 8'd120}: color_data = 12'h06b;
			{8'd66, 8'd121}: color_data = 12'h06b;
			{8'd66, 8'd122}: color_data = 12'h06b;
			{8'd66, 8'd123}: color_data = 12'h06b;
			{8'd66, 8'd124}: color_data = 12'h06b;
			{8'd66, 8'd125}: color_data = 12'h06b;
			{8'd66, 8'd126}: color_data = 12'h05a;
			{8'd66, 8'd127}: color_data = 12'h047;
			{8'd66, 8'd128}: color_data = 12'h234;
			{8'd66, 8'd129}: color_data = 12'h433;
			{8'd66, 8'd130}: color_data = 12'h531;
			{8'd66, 8'd131}: color_data = 12'h521;
			{8'd66, 8'd132}: color_data = 12'h321;
			{8'd66, 8'd133}: color_data = 12'h000;
			{8'd67, 8'd14}: color_data = 12'hfc6;
			{8'd67, 8'd15}: color_data = 12'hfc5;
			{8'd67, 8'd16}: color_data = 12'hfc5;
			{8'd67, 8'd17}: color_data = 12'hfc5;
			{8'd67, 8'd18}: color_data = 12'heb2;
			{8'd67, 8'd19}: color_data = 12'hd90;
			{8'd67, 8'd20}: color_data = 12'hd90;
			{8'd67, 8'd21}: color_data = 12'hd90;
			{8'd67, 8'd22}: color_data = 12'hd90;
			{8'd67, 8'd23}: color_data = 12'hd90;
			{8'd67, 8'd24}: color_data = 12'hd90;
			{8'd67, 8'd25}: color_data = 12'hd90;
			{8'd67, 8'd26}: color_data = 12'hea1;
			{8'd67, 8'd27}: color_data = 12'hfc5;
			{8'd67, 8'd28}: color_data = 12'hfc5;
			{8'd67, 8'd29}: color_data = 12'hfd6;
			{8'd67, 8'd57}: color_data = 12'h500;
			{8'd67, 8'd58}: color_data = 12'hd12;
			{8'd67, 8'd59}: color_data = 12'he12;
			{8'd67, 8'd60}: color_data = 12'he12;
			{8'd67, 8'd61}: color_data = 12'hc12;
			{8'd67, 8'd62}: color_data = 12'h911;
			{8'd67, 8'd63}: color_data = 12'h400;
			{8'd67, 8'd64}: color_data = 12'h000;
			{8'd67, 8'd89}: color_data = 12'h300;
			{8'd67, 8'd90}: color_data = 12'ha12;
			{8'd67, 8'd91}: color_data = 12'ha33;
			{8'd67, 8'd92}: color_data = 12'h945;
			{8'd67, 8'd93}: color_data = 12'h956;
			{8'd67, 8'd94}: color_data = 12'h956;
			{8'd67, 8'd95}: color_data = 12'h955;
			{8'd67, 8'd96}: color_data = 12'ha23;
			{8'd67, 8'd97}: color_data = 12'hc11;
			{8'd67, 8'd98}: color_data = 12'hf12;
			{8'd67, 8'd99}: color_data = 12'hf12;
			{8'd67, 8'd100}: color_data = 12'h911;
			{8'd67, 8'd101}: color_data = 12'h000;
			{8'd67, 8'd106}: color_data = 12'h000;
			{8'd67, 8'd107}: color_data = 12'h036;
			{8'd67, 8'd108}: color_data = 12'h06b;
			{8'd67, 8'd109}: color_data = 12'h06b;
			{8'd67, 8'd110}: color_data = 12'h06b;
			{8'd67, 8'd111}: color_data = 12'h06b;
			{8'd67, 8'd112}: color_data = 12'h06b;
			{8'd67, 8'd113}: color_data = 12'h06b;
			{8'd67, 8'd114}: color_data = 12'h06b;
			{8'd67, 8'd115}: color_data = 12'h06b;
			{8'd67, 8'd116}: color_data = 12'h06b;
			{8'd67, 8'd117}: color_data = 12'h06b;
			{8'd67, 8'd118}: color_data = 12'h06b;
			{8'd67, 8'd119}: color_data = 12'h06b;
			{8'd67, 8'd120}: color_data = 12'h06b;
			{8'd67, 8'd121}: color_data = 12'h06b;
			{8'd67, 8'd122}: color_data = 12'h06b;
			{8'd67, 8'd123}: color_data = 12'h06b;
			{8'd67, 8'd124}: color_data = 12'h06b;
			{8'd67, 8'd125}: color_data = 12'h06b;
			{8'd67, 8'd126}: color_data = 12'h06b;
			{8'd67, 8'd127}: color_data = 12'h06b;
			{8'd67, 8'd128}: color_data = 12'h06a;
			{8'd67, 8'd129}: color_data = 12'h036;
			{8'd67, 8'd130}: color_data = 12'h000;
			{8'd67, 8'd131}: color_data = 12'h000;
			{8'd68, 8'd14}: color_data = 12'hfc5;
			{8'd68, 8'd15}: color_data = 12'hfc5;
			{8'd68, 8'd16}: color_data = 12'hfc4;
			{8'd68, 8'd17}: color_data = 12'hea0;
			{8'd68, 8'd18}: color_data = 12'hd90;
			{8'd68, 8'd19}: color_data = 12'hd90;
			{8'd68, 8'd20}: color_data = 12'hd90;
			{8'd68, 8'd21}: color_data = 12'hd90;
			{8'd68, 8'd22}: color_data = 12'hd90;
			{8'd68, 8'd23}: color_data = 12'hd90;
			{8'd68, 8'd24}: color_data = 12'hea1;
			{8'd68, 8'd25}: color_data = 12'heb2;
			{8'd68, 8'd26}: color_data = 12'hfb3;
			{8'd68, 8'd27}: color_data = 12'hfc5;
			{8'd68, 8'd28}: color_data = 12'hfc4;
			{8'd68, 8'd56}: color_data = 12'h000;
			{8'd68, 8'd57}: color_data = 12'hb11;
			{8'd68, 8'd58}: color_data = 12'hf12;
			{8'd68, 8'd59}: color_data = 12'he12;
			{8'd68, 8'd60}: color_data = 12'he12;
			{8'd68, 8'd61}: color_data = 12'hf12;
			{8'd68, 8'd62}: color_data = 12'hf12;
			{8'd68, 8'd63}: color_data = 12'he12;
			{8'd68, 8'd64}: color_data = 12'h801;
			{8'd68, 8'd65}: color_data = 12'h100;
			{8'd68, 8'd88}: color_data = 12'h222;
			{8'd68, 8'd89}: color_data = 12'h988;
			{8'd68, 8'd90}: color_data = 12'hddd;
			{8'd68, 8'd91}: color_data = 12'hfff;
			{8'd68, 8'd92}: color_data = 12'hfff;
			{8'd68, 8'd93}: color_data = 12'hfff;
			{8'd68, 8'd94}: color_data = 12'hfff;
			{8'd68, 8'd95}: color_data = 12'hfff;
			{8'd68, 8'd96}: color_data = 12'heff;
			{8'd68, 8'd97}: color_data = 12'ha88;
			{8'd68, 8'd98}: color_data = 12'hb11;
			{8'd68, 8'd99}: color_data = 12'hf12;
			{8'd68, 8'd100}: color_data = 12'hb11;
			{8'd68, 8'd101}: color_data = 12'h000;
			{8'd68, 8'd105}: color_data = 12'h000;
			{8'd68, 8'd106}: color_data = 12'h000;
			{8'd68, 8'd107}: color_data = 12'h012;
			{8'd68, 8'd108}: color_data = 12'h05a;
			{8'd68, 8'd109}: color_data = 12'h06b;
			{8'd68, 8'd110}: color_data = 12'h06b;
			{8'd68, 8'd111}: color_data = 12'h06b;
			{8'd68, 8'd112}: color_data = 12'h06b;
			{8'd68, 8'd113}: color_data = 12'h06b;
			{8'd68, 8'd114}: color_data = 12'h06b;
			{8'd68, 8'd115}: color_data = 12'h06b;
			{8'd68, 8'd116}: color_data = 12'h06b;
			{8'd68, 8'd117}: color_data = 12'h06b;
			{8'd68, 8'd118}: color_data = 12'h06b;
			{8'd68, 8'd119}: color_data = 12'h06b;
			{8'd68, 8'd120}: color_data = 12'h06b;
			{8'd68, 8'd121}: color_data = 12'h06a;
			{8'd68, 8'd122}: color_data = 12'h059;
			{8'd68, 8'd123}: color_data = 12'h047;
			{8'd68, 8'd124}: color_data = 12'h036;
			{8'd68, 8'd125}: color_data = 12'h036;
			{8'd68, 8'd126}: color_data = 12'h025;
			{8'd68, 8'd127}: color_data = 12'h024;
			{8'd68, 8'd128}: color_data = 12'h012;
			{8'd68, 8'd129}: color_data = 12'h000;
			{8'd69, 8'd14}: color_data = 12'hfc5;
			{8'd69, 8'd15}: color_data = 12'hfc5;
			{8'd69, 8'd16}: color_data = 12'hfb3;
			{8'd69, 8'd17}: color_data = 12'hd90;
			{8'd69, 8'd18}: color_data = 12'hd90;
			{8'd69, 8'd19}: color_data = 12'hd90;
			{8'd69, 8'd20}: color_data = 12'hd90;
			{8'd69, 8'd21}: color_data = 12'hd90;
			{8'd69, 8'd22}: color_data = 12'hd90;
			{8'd69, 8'd23}: color_data = 12'hfb3;
			{8'd69, 8'd24}: color_data = 12'hfc6;
			{8'd69, 8'd25}: color_data = 12'hfc6;
			{8'd69, 8'd26}: color_data = 12'hfc5;
			{8'd69, 8'd27}: color_data = 12'hfc5;
			{8'd69, 8'd28}: color_data = 12'hfc5;
			{8'd69, 8'd56}: color_data = 12'h300;
			{8'd69, 8'd57}: color_data = 12'hd12;
			{8'd69, 8'd58}: color_data = 12'hf12;
			{8'd69, 8'd59}: color_data = 12'he12;
			{8'd69, 8'd60}: color_data = 12'he12;
			{8'd69, 8'd61}: color_data = 12'he12;
			{8'd69, 8'd62}: color_data = 12'he12;
			{8'd69, 8'd63}: color_data = 12'hf12;
			{8'd69, 8'd64}: color_data = 12'hf12;
			{8'd69, 8'd65}: color_data = 12'h911;
			{8'd69, 8'd66}: color_data = 12'h000;
			{8'd69, 8'd87}: color_data = 12'h222;
			{8'd69, 8'd88}: color_data = 12'hccc;
			{8'd69, 8'd89}: color_data = 12'hfff;
			{8'd69, 8'd90}: color_data = 12'hccc;
			{8'd69, 8'd91}: color_data = 12'hbbb;
			{8'd69, 8'd92}: color_data = 12'hbbb;
			{8'd69, 8'd93}: color_data = 12'hddd;
			{8'd69, 8'd94}: color_data = 12'hfff;
			{8'd69, 8'd95}: color_data = 12'hfff;
			{8'd69, 8'd96}: color_data = 12'hfff;
			{8'd69, 8'd97}: color_data = 12'hfff;
			{8'd69, 8'd98}: color_data = 12'h977;
			{8'd69, 8'd99}: color_data = 12'hd01;
			{8'd69, 8'd100}: color_data = 12'hd11;
			{8'd69, 8'd101}: color_data = 12'h200;
			{8'd69, 8'd102}: color_data = 12'h000;
			{8'd69, 8'd103}: color_data = 12'h012;
			{8'd69, 8'd104}: color_data = 12'h024;
			{8'd69, 8'd105}: color_data = 12'h035;
			{8'd69, 8'd106}: color_data = 12'h047;
			{8'd69, 8'd107}: color_data = 12'h047;
			{8'd69, 8'd108}: color_data = 12'h047;
			{8'd69, 8'd109}: color_data = 12'h06b;
			{8'd69, 8'd110}: color_data = 12'h06b;
			{8'd69, 8'd111}: color_data = 12'h06b;
			{8'd69, 8'd112}: color_data = 12'h06b;
			{8'd69, 8'd113}: color_data = 12'h06b;
			{8'd69, 8'd114}: color_data = 12'h06b;
			{8'd69, 8'd115}: color_data = 12'h06b;
			{8'd69, 8'd116}: color_data = 12'h06b;
			{8'd69, 8'd117}: color_data = 12'h06b;
			{8'd69, 8'd118}: color_data = 12'h06b;
			{8'd69, 8'd119}: color_data = 12'h05a;
			{8'd69, 8'd120}: color_data = 12'h036;
			{8'd69, 8'd121}: color_data = 12'h013;
			{8'd69, 8'd122}: color_data = 12'h000;
			{8'd69, 8'd123}: color_data = 12'h000;
			{8'd69, 8'd124}: color_data = 12'h000;
			{8'd70, 8'd12}: color_data = 12'hff0;
			{8'd70, 8'd13}: color_data = 12'hfd6;
			{8'd70, 8'd14}: color_data = 12'hfc6;
			{8'd70, 8'd15}: color_data = 12'hfc5;
			{8'd70, 8'd16}: color_data = 12'hfc5;
			{8'd70, 8'd17}: color_data = 12'hfb3;
			{8'd70, 8'd18}: color_data = 12'hd90;
			{8'd70, 8'd19}: color_data = 12'hd90;
			{8'd70, 8'd20}: color_data = 12'hd90;
			{8'd70, 8'd21}: color_data = 12'hd90;
			{8'd70, 8'd22}: color_data = 12'hd90;
			{8'd70, 8'd23}: color_data = 12'hda0;
			{8'd70, 8'd24}: color_data = 12'heb2;
			{8'd70, 8'd25}: color_data = 12'hfc4;
			{8'd70, 8'd26}: color_data = 12'hfc5;
			{8'd70, 8'd27}: color_data = 12'hfc5;
			{8'd70, 8'd56}: color_data = 12'h400;
			{8'd70, 8'd57}: color_data = 12'he12;
			{8'd70, 8'd58}: color_data = 12'hf12;
			{8'd70, 8'd59}: color_data = 12'he12;
			{8'd70, 8'd60}: color_data = 12'he12;
			{8'd70, 8'd61}: color_data = 12'he12;
			{8'd70, 8'd62}: color_data = 12'he12;
			{8'd70, 8'd63}: color_data = 12'he12;
			{8'd70, 8'd64}: color_data = 12'he12;
			{8'd70, 8'd65}: color_data = 12'hf12;
			{8'd70, 8'd66}: color_data = 12'h801;
			{8'd70, 8'd67}: color_data = 12'h000;
			{8'd70, 8'd85}: color_data = 12'h000;
			{8'd70, 8'd86}: color_data = 12'h000;
			{8'd70, 8'd87}: color_data = 12'h555;
			{8'd70, 8'd88}: color_data = 12'hbbb;
			{8'd70, 8'd89}: color_data = 12'h999;
			{8'd70, 8'd90}: color_data = 12'hccc;
			{8'd70, 8'd91}: color_data = 12'hddd;
			{8'd70, 8'd92}: color_data = 12'hddd;
			{8'd70, 8'd93}: color_data = 12'heee;
			{8'd70, 8'd94}: color_data = 12'hfff;
			{8'd70, 8'd95}: color_data = 12'hfff;
			{8'd70, 8'd96}: color_data = 12'hbbb;
			{8'd70, 8'd97}: color_data = 12'h987;
			{8'd70, 8'd98}: color_data = 12'h876;
			{8'd70, 8'd99}: color_data = 12'h632;
			{8'd70, 8'd100}: color_data = 12'h223;
			{8'd70, 8'd101}: color_data = 12'h036;
			{8'd70, 8'd102}: color_data = 12'h048;
			{8'd70, 8'd103}: color_data = 12'h05a;
			{8'd70, 8'd104}: color_data = 12'h06b;
			{8'd70, 8'd105}: color_data = 12'h06b;
			{8'd70, 8'd106}: color_data = 12'h06b;
			{8'd70, 8'd107}: color_data = 12'h06b;
			{8'd70, 8'd108}: color_data = 12'h047;
			{8'd70, 8'd109}: color_data = 12'h059;
			{8'd70, 8'd110}: color_data = 12'h06b;
			{8'd70, 8'd111}: color_data = 12'h06b;
			{8'd70, 8'd112}: color_data = 12'h06b;
			{8'd70, 8'd113}: color_data = 12'h06b;
			{8'd70, 8'd114}: color_data = 12'h06b;
			{8'd70, 8'd115}: color_data = 12'h06b;
			{8'd70, 8'd116}: color_data = 12'h06b;
			{8'd70, 8'd117}: color_data = 12'h06b;
			{8'd70, 8'd118}: color_data = 12'h059;
			{8'd70, 8'd119}: color_data = 12'h012;
			{8'd70, 8'd120}: color_data = 12'h000;
			{8'd71, 8'd10}: color_data = 12'hfc5;
			{8'd71, 8'd11}: color_data = 12'hfc5;
			{8'd71, 8'd12}: color_data = 12'hfc5;
			{8'd71, 8'd13}: color_data = 12'hfc5;
			{8'd71, 8'd14}: color_data = 12'hfc5;
			{8'd71, 8'd15}: color_data = 12'hfc5;
			{8'd71, 8'd16}: color_data = 12'hfc5;
			{8'd71, 8'd17}: color_data = 12'hfc6;
			{8'd71, 8'd18}: color_data = 12'heb2;
			{8'd71, 8'd19}: color_data = 12'hd90;
			{8'd71, 8'd20}: color_data = 12'hd90;
			{8'd71, 8'd21}: color_data = 12'hd90;
			{8'd71, 8'd22}: color_data = 12'hd90;
			{8'd71, 8'd23}: color_data = 12'hd90;
			{8'd71, 8'd24}: color_data = 12'hd90;
			{8'd71, 8'd25}: color_data = 12'hea1;
			{8'd71, 8'd26}: color_data = 12'hfc5;
			{8'd71, 8'd27}: color_data = 12'hfc5;
			{8'd71, 8'd28}: color_data = 12'hfb5;
			{8'd71, 8'd56}: color_data = 12'h400;
			{8'd71, 8'd57}: color_data = 12'he12;
			{8'd71, 8'd58}: color_data = 12'hf12;
			{8'd71, 8'd59}: color_data = 12'he12;
			{8'd71, 8'd60}: color_data = 12'he12;
			{8'd71, 8'd61}: color_data = 12'he12;
			{8'd71, 8'd62}: color_data = 12'he12;
			{8'd71, 8'd63}: color_data = 12'he12;
			{8'd71, 8'd64}: color_data = 12'he12;
			{8'd71, 8'd65}: color_data = 12'hf12;
			{8'd71, 8'd66}: color_data = 12'hd12;
			{8'd71, 8'd67}: color_data = 12'h200;
			{8'd71, 8'd84}: color_data = 12'h000;
			{8'd71, 8'd85}: color_data = 12'h555;
			{8'd71, 8'd86}: color_data = 12'hccc;
			{8'd71, 8'd87}: color_data = 12'heee;
			{8'd71, 8'd88}: color_data = 12'hfff;
			{8'd71, 8'd89}: color_data = 12'hfff;
			{8'd71, 8'd90}: color_data = 12'hfff;
			{8'd71, 8'd91}: color_data = 12'hfff;
			{8'd71, 8'd92}: color_data = 12'hfff;
			{8'd71, 8'd93}: color_data = 12'hfff;
			{8'd71, 8'd94}: color_data = 12'hbbb;
			{8'd71, 8'd95}: color_data = 12'h876;
			{8'd71, 8'd96}: color_data = 12'ha76;
			{8'd71, 8'd97}: color_data = 12'hc97;
			{8'd71, 8'd98}: color_data = 12'h965;
			{8'd71, 8'd99}: color_data = 12'h147;
			{8'd71, 8'd100}: color_data = 12'h06b;
			{8'd71, 8'd101}: color_data = 12'h06b;
			{8'd71, 8'd102}: color_data = 12'h06b;
			{8'd71, 8'd103}: color_data = 12'h06b;
			{8'd71, 8'd104}: color_data = 12'h06b;
			{8'd71, 8'd105}: color_data = 12'h06b;
			{8'd71, 8'd106}: color_data = 12'h06b;
			{8'd71, 8'd107}: color_data = 12'h06b;
			{8'd71, 8'd108}: color_data = 12'h05a;
			{8'd71, 8'd109}: color_data = 12'h047;
			{8'd71, 8'd110}: color_data = 12'h06b;
			{8'd71, 8'd111}: color_data = 12'h06b;
			{8'd71, 8'd112}: color_data = 12'h06b;
			{8'd71, 8'd113}: color_data = 12'h06b;
			{8'd71, 8'd114}: color_data = 12'h06b;
			{8'd71, 8'd115}: color_data = 12'h06b;
			{8'd71, 8'd116}: color_data = 12'h06b;
			{8'd71, 8'd117}: color_data = 12'h06b;
			{8'd71, 8'd118}: color_data = 12'h059;
			{8'd71, 8'd119}: color_data = 12'h001;
			{8'd72, 8'd9}: color_data = 12'hfc4;
			{8'd72, 8'd10}: color_data = 12'hfc4;
			{8'd72, 8'd11}: color_data = 12'hfc5;
			{8'd72, 8'd12}: color_data = 12'hfc5;
			{8'd72, 8'd13}: color_data = 12'hfc4;
			{8'd72, 8'd14}: color_data = 12'hfc4;
			{8'd72, 8'd15}: color_data = 12'hfb3;
			{8'd72, 8'd16}: color_data = 12'heb2;
			{8'd72, 8'd17}: color_data = 12'hea1;
			{8'd72, 8'd18}: color_data = 12'hea0;
			{8'd72, 8'd19}: color_data = 12'hd90;
			{8'd72, 8'd20}: color_data = 12'hd90;
			{8'd72, 8'd21}: color_data = 12'hd90;
			{8'd72, 8'd22}: color_data = 12'hd90;
			{8'd72, 8'd23}: color_data = 12'hd90;
			{8'd72, 8'd24}: color_data = 12'hd90;
			{8'd72, 8'd25}: color_data = 12'hea1;
			{8'd72, 8'd26}: color_data = 12'hfc5;
			{8'd72, 8'd27}: color_data = 12'hfc5;
			{8'd72, 8'd28}: color_data = 12'hff5;
			{8'd72, 8'd56}: color_data = 12'h400;
			{8'd72, 8'd57}: color_data = 12'he12;
			{8'd72, 8'd58}: color_data = 12'hf12;
			{8'd72, 8'd59}: color_data = 12'he12;
			{8'd72, 8'd60}: color_data = 12'he12;
			{8'd72, 8'd61}: color_data = 12'he12;
			{8'd72, 8'd62}: color_data = 12'he12;
			{8'd72, 8'd63}: color_data = 12'he12;
			{8'd72, 8'd64}: color_data = 12'he12;
			{8'd72, 8'd65}: color_data = 12'he12;
			{8'd72, 8'd66}: color_data = 12'hf12;
			{8'd72, 8'd67}: color_data = 12'h601;
			{8'd72, 8'd82}: color_data = 12'h000;
			{8'd72, 8'd83}: color_data = 12'h000;
			{8'd72, 8'd84}: color_data = 12'h555;
			{8'd72, 8'd85}: color_data = 12'heee;
			{8'd72, 8'd86}: color_data = 12'hfff;
			{8'd72, 8'd87}: color_data = 12'hfff;
			{8'd72, 8'd88}: color_data = 12'hfff;
			{8'd72, 8'd89}: color_data = 12'hfff;
			{8'd72, 8'd90}: color_data = 12'hfff;
			{8'd72, 8'd91}: color_data = 12'hfff;
			{8'd72, 8'd92}: color_data = 12'hfff;
			{8'd72, 8'd93}: color_data = 12'h877;
			{8'd72, 8'd94}: color_data = 12'h975;
			{8'd72, 8'd95}: color_data = 12'hc97;
			{8'd72, 8'd96}: color_data = 12'hc97;
			{8'd72, 8'd97}: color_data = 12'h555;
			{8'd72, 8'd98}: color_data = 12'h048;
			{8'd72, 8'd99}: color_data = 12'h06b;
			{8'd72, 8'd100}: color_data = 12'h06b;
			{8'd72, 8'd101}: color_data = 12'h06b;
			{8'd72, 8'd102}: color_data = 12'h06b;
			{8'd72, 8'd103}: color_data = 12'h06b;
			{8'd72, 8'd104}: color_data = 12'h06b;
			{8'd72, 8'd105}: color_data = 12'h06b;
			{8'd72, 8'd106}: color_data = 12'h06b;
			{8'd72, 8'd107}: color_data = 12'h06b;
			{8'd72, 8'd108}: color_data = 12'h06b;
			{8'd72, 8'd109}: color_data = 12'h058;
			{8'd72, 8'd110}: color_data = 12'h06a;
			{8'd72, 8'd111}: color_data = 12'h06b;
			{8'd72, 8'd112}: color_data = 12'h06b;
			{8'd72, 8'd113}: color_data = 12'h06b;
			{8'd72, 8'd114}: color_data = 12'h06b;
			{8'd72, 8'd115}: color_data = 12'h06b;
			{8'd72, 8'd116}: color_data = 12'h06b;
			{8'd72, 8'd117}: color_data = 12'h06b;
			{8'd72, 8'd118}: color_data = 12'h06a;
			{8'd72, 8'd119}: color_data = 12'h013;
			{8'd73, 8'd9}: color_data = 12'hfc4;
			{8'd73, 8'd10}: color_data = 12'hfc5;
			{8'd73, 8'd11}: color_data = 12'hfc4;
			{8'd73, 8'd12}: color_data = 12'hea1;
			{8'd73, 8'd13}: color_data = 12'hda0;
			{8'd73, 8'd14}: color_data = 12'hd90;
			{8'd73, 8'd15}: color_data = 12'hd90;
			{8'd73, 8'd16}: color_data = 12'hd90;
			{8'd73, 8'd17}: color_data = 12'hd90;
			{8'd73, 8'd18}: color_data = 12'hd90;
			{8'd73, 8'd19}: color_data = 12'hd90;
			{8'd73, 8'd20}: color_data = 12'hd90;
			{8'd73, 8'd21}: color_data = 12'hd90;
			{8'd73, 8'd22}: color_data = 12'hd90;
			{8'd73, 8'd23}: color_data = 12'hd90;
			{8'd73, 8'd24}: color_data = 12'hd90;
			{8'd73, 8'd25}: color_data = 12'heb2;
			{8'd73, 8'd26}: color_data = 12'hfc5;
			{8'd73, 8'd27}: color_data = 12'hfc5;
			{8'd73, 8'd56}: color_data = 12'h300;
			{8'd73, 8'd57}: color_data = 12'hd12;
			{8'd73, 8'd58}: color_data = 12'hf12;
			{8'd73, 8'd59}: color_data = 12'he12;
			{8'd73, 8'd60}: color_data = 12'he12;
			{8'd73, 8'd61}: color_data = 12'he12;
			{8'd73, 8'd62}: color_data = 12'he12;
			{8'd73, 8'd63}: color_data = 12'he12;
			{8'd73, 8'd64}: color_data = 12'he12;
			{8'd73, 8'd65}: color_data = 12'he12;
			{8'd73, 8'd66}: color_data = 12'hf12;
			{8'd73, 8'd67}: color_data = 12'h811;
			{8'd73, 8'd68}: color_data = 12'h000;
			{8'd73, 8'd81}: color_data = 12'h222;
			{8'd73, 8'd82}: color_data = 12'h888;
			{8'd73, 8'd83}: color_data = 12'hccc;
			{8'd73, 8'd84}: color_data = 12'heee;
			{8'd73, 8'd85}: color_data = 12'hfff;
			{8'd73, 8'd86}: color_data = 12'hfff;
			{8'd73, 8'd87}: color_data = 12'hfff;
			{8'd73, 8'd88}: color_data = 12'hfff;
			{8'd73, 8'd89}: color_data = 12'hfff;
			{8'd73, 8'd90}: color_data = 12'hfff;
			{8'd73, 8'd91}: color_data = 12'hfff;
			{8'd73, 8'd92}: color_data = 12'hfff;
			{8'd73, 8'd93}: color_data = 12'h877;
			{8'd73, 8'd94}: color_data = 12'hd97;
			{8'd73, 8'd95}: color_data = 12'ha76;
			{8'd73, 8'd96}: color_data = 12'h345;
			{8'd73, 8'd97}: color_data = 12'h05a;
			{8'd73, 8'd98}: color_data = 12'h06b;
			{8'd73, 8'd99}: color_data = 12'h06b;
			{8'd73, 8'd100}: color_data = 12'h06b;
			{8'd73, 8'd101}: color_data = 12'h06b;
			{8'd73, 8'd102}: color_data = 12'h06b;
			{8'd73, 8'd103}: color_data = 12'h06b;
			{8'd73, 8'd104}: color_data = 12'h06b;
			{8'd73, 8'd105}: color_data = 12'h06b;
			{8'd73, 8'd106}: color_data = 12'h06b;
			{8'd73, 8'd107}: color_data = 12'h06b;
			{8'd73, 8'd108}: color_data = 12'h06b;
			{8'd73, 8'd109}: color_data = 12'h06b;
			{8'd73, 8'd110}: color_data = 12'h06b;
			{8'd73, 8'd111}: color_data = 12'h06b;
			{8'd73, 8'd112}: color_data = 12'h06b;
			{8'd73, 8'd113}: color_data = 12'h06b;
			{8'd73, 8'd114}: color_data = 12'h06b;
			{8'd73, 8'd115}: color_data = 12'h06b;
			{8'd73, 8'd116}: color_data = 12'h06b;
			{8'd73, 8'd117}: color_data = 12'h06b;
			{8'd73, 8'd118}: color_data = 12'h06b;
			{8'd73, 8'd119}: color_data = 12'h024;
			{8'd74, 8'd9}: color_data = 12'hfc5;
			{8'd74, 8'd10}: color_data = 12'hfc5;
			{8'd74, 8'd11}: color_data = 12'hfc4;
			{8'd74, 8'd12}: color_data = 12'hd90;
			{8'd74, 8'd13}: color_data = 12'hd90;
			{8'd74, 8'd14}: color_data = 12'hd90;
			{8'd74, 8'd15}: color_data = 12'hd90;
			{8'd74, 8'd16}: color_data = 12'hd90;
			{8'd74, 8'd17}: color_data = 12'hd90;
			{8'd74, 8'd18}: color_data = 12'hd90;
			{8'd74, 8'd19}: color_data = 12'hd90;
			{8'd74, 8'd20}: color_data = 12'hd90;
			{8'd74, 8'd21}: color_data = 12'hd90;
			{8'd74, 8'd22}: color_data = 12'hd90;
			{8'd74, 8'd23}: color_data = 12'hd90;
			{8'd74, 8'd24}: color_data = 12'hea0;
			{8'd74, 8'd25}: color_data = 12'hfc4;
			{8'd74, 8'd26}: color_data = 12'hfc4;
			{8'd74, 8'd27}: color_data = 12'hfc4;
			{8'd74, 8'd56}: color_data = 12'h200;
			{8'd74, 8'd57}: color_data = 12'hc12;
			{8'd74, 8'd58}: color_data = 12'hf12;
			{8'd74, 8'd59}: color_data = 12'he12;
			{8'd74, 8'd60}: color_data = 12'he12;
			{8'd74, 8'd61}: color_data = 12'he12;
			{8'd74, 8'd62}: color_data = 12'he12;
			{8'd74, 8'd63}: color_data = 12'he12;
			{8'd74, 8'd64}: color_data = 12'he12;
			{8'd74, 8'd65}: color_data = 12'he12;
			{8'd74, 8'd66}: color_data = 12'hf12;
			{8'd74, 8'd67}: color_data = 12'ha11;
			{8'd74, 8'd68}: color_data = 12'h000;
			{8'd74, 8'd80}: color_data = 12'h111;
			{8'd74, 8'd81}: color_data = 12'hbbb;
			{8'd74, 8'd82}: color_data = 12'hfff;
			{8'd74, 8'd83}: color_data = 12'hfff;
			{8'd74, 8'd84}: color_data = 12'hfff;
			{8'd74, 8'd85}: color_data = 12'hfff;
			{8'd74, 8'd86}: color_data = 12'hfff;
			{8'd74, 8'd87}: color_data = 12'hddd;
			{8'd74, 8'd88}: color_data = 12'hfff;
			{8'd74, 8'd89}: color_data = 12'hccc;
			{8'd74, 8'd90}: color_data = 12'hddd;
			{8'd74, 8'd91}: color_data = 12'hfff;
			{8'd74, 8'd92}: color_data = 12'hfff;
			{8'd74, 8'd93}: color_data = 12'ha99;
			{8'd74, 8'd94}: color_data = 12'h754;
			{8'd74, 8'd95}: color_data = 12'h147;
			{8'd74, 8'd96}: color_data = 12'h06b;
			{8'd74, 8'd97}: color_data = 12'h06b;
			{8'd74, 8'd98}: color_data = 12'h06b;
			{8'd74, 8'd99}: color_data = 12'h06b;
			{8'd74, 8'd100}: color_data = 12'h06b;
			{8'd74, 8'd101}: color_data = 12'h06b;
			{8'd74, 8'd102}: color_data = 12'h06b;
			{8'd74, 8'd103}: color_data = 12'h06b;
			{8'd74, 8'd104}: color_data = 12'h06b;
			{8'd74, 8'd105}: color_data = 12'h06b;
			{8'd74, 8'd106}: color_data = 12'h06b;
			{8'd74, 8'd107}: color_data = 12'h06b;
			{8'd74, 8'd108}: color_data = 12'h06b;
			{8'd74, 8'd109}: color_data = 12'h06b;
			{8'd74, 8'd110}: color_data = 12'h06b;
			{8'd74, 8'd111}: color_data = 12'h06b;
			{8'd74, 8'd112}: color_data = 12'h06b;
			{8'd74, 8'd113}: color_data = 12'h06b;
			{8'd74, 8'd114}: color_data = 12'h06b;
			{8'd74, 8'd115}: color_data = 12'h06b;
			{8'd74, 8'd116}: color_data = 12'h06b;
			{8'd74, 8'd117}: color_data = 12'h06b;
			{8'd74, 8'd118}: color_data = 12'h06b;
			{8'd74, 8'd119}: color_data = 12'h035;
			{8'd75, 8'd9}: color_data = 12'hfc5;
			{8'd75, 8'd10}: color_data = 12'hfc5;
			{8'd75, 8'd11}: color_data = 12'hfc4;
			{8'd75, 8'd12}: color_data = 12'hd90;
			{8'd75, 8'd13}: color_data = 12'hd90;
			{8'd75, 8'd14}: color_data = 12'hd90;
			{8'd75, 8'd15}: color_data = 12'hd90;
			{8'd75, 8'd16}: color_data = 12'hd90;
			{8'd75, 8'd17}: color_data = 12'hd90;
			{8'd75, 8'd18}: color_data = 12'hd90;
			{8'd75, 8'd19}: color_data = 12'hd90;
			{8'd75, 8'd20}: color_data = 12'hea0;
			{8'd75, 8'd21}: color_data = 12'hea1;
			{8'd75, 8'd22}: color_data = 12'heb2;
			{8'd75, 8'd23}: color_data = 12'hfb3;
			{8'd75, 8'd24}: color_data = 12'hfc5;
			{8'd75, 8'd25}: color_data = 12'hfc5;
			{8'd75, 8'd26}: color_data = 12'hfc4;
			{8'd75, 8'd27}: color_data = 12'hfc5;
			{8'd75, 8'd56}: color_data = 12'h000;
			{8'd75, 8'd57}: color_data = 12'hb11;
			{8'd75, 8'd58}: color_data = 12'he12;
			{8'd75, 8'd59}: color_data = 12'he12;
			{8'd75, 8'd60}: color_data = 12'he12;
			{8'd75, 8'd61}: color_data = 12'he12;
			{8'd75, 8'd62}: color_data = 12'he12;
			{8'd75, 8'd63}: color_data = 12'he12;
			{8'd75, 8'd64}: color_data = 12'he12;
			{8'd75, 8'd65}: color_data = 12'he12;
			{8'd75, 8'd66}: color_data = 12'hf12;
			{8'd75, 8'd67}: color_data = 12'ha11;
			{8'd75, 8'd68}: color_data = 12'h000;
			{8'd75, 8'd80}: color_data = 12'h666;
			{8'd75, 8'd81}: color_data = 12'hfff;
			{8'd75, 8'd82}: color_data = 12'hfff;
			{8'd75, 8'd83}: color_data = 12'hfff;
			{8'd75, 8'd84}: color_data = 12'hfff;
			{8'd75, 8'd85}: color_data = 12'hfff;
			{8'd75, 8'd86}: color_data = 12'hfff;
			{8'd75, 8'd87}: color_data = 12'haaa;
			{8'd75, 8'd88}: color_data = 12'hfff;
			{8'd75, 8'd89}: color_data = 12'hddd;
			{8'd75, 8'd90}: color_data = 12'hbbb;
			{8'd75, 8'd91}: color_data = 12'hfff;
			{8'd75, 8'd92}: color_data = 12'hfff;
			{8'd75, 8'd93}: color_data = 12'haaa;
			{8'd75, 8'd94}: color_data = 12'h047;
			{8'd75, 8'd95}: color_data = 12'h06b;
			{8'd75, 8'd96}: color_data = 12'h06a;
			{8'd75, 8'd97}: color_data = 12'h06b;
			{8'd75, 8'd98}: color_data = 12'h06b;
			{8'd75, 8'd99}: color_data = 12'h06b;
			{8'd75, 8'd100}: color_data = 12'h06b;
			{8'd75, 8'd101}: color_data = 12'h06b;
			{8'd75, 8'd102}: color_data = 12'h06b;
			{8'd75, 8'd103}: color_data = 12'h06b;
			{8'd75, 8'd104}: color_data = 12'h06b;
			{8'd75, 8'd105}: color_data = 12'h06b;
			{8'd75, 8'd106}: color_data = 12'h06b;
			{8'd75, 8'd107}: color_data = 12'h06b;
			{8'd75, 8'd108}: color_data = 12'h06b;
			{8'd75, 8'd109}: color_data = 12'h06b;
			{8'd75, 8'd110}: color_data = 12'h06b;
			{8'd75, 8'd111}: color_data = 12'h06b;
			{8'd75, 8'd112}: color_data = 12'h06b;
			{8'd75, 8'd113}: color_data = 12'h06b;
			{8'd75, 8'd114}: color_data = 12'h06b;
			{8'd75, 8'd115}: color_data = 12'h06b;
			{8'd75, 8'd116}: color_data = 12'h06b;
			{8'd75, 8'd117}: color_data = 12'h06b;
			{8'd75, 8'd118}: color_data = 12'h06b;
			{8'd75, 8'd119}: color_data = 12'h036;
			{8'd75, 8'd120}: color_data = 12'h000;
			{8'd76, 8'd9}: color_data = 12'hfc5;
			{8'd76, 8'd10}: color_data = 12'hfc5;
			{8'd76, 8'd11}: color_data = 12'hfc4;
			{8'd76, 8'd12}: color_data = 12'hd90;
			{8'd76, 8'd13}: color_data = 12'hd90;
			{8'd76, 8'd14}: color_data = 12'hd90;
			{8'd76, 8'd15}: color_data = 12'hd90;
			{8'd76, 8'd16}: color_data = 12'hda0;
			{8'd76, 8'd17}: color_data = 12'hea1;
			{8'd76, 8'd18}: color_data = 12'heb2;
			{8'd76, 8'd19}: color_data = 12'hfb3;
			{8'd76, 8'd20}: color_data = 12'hfc4;
			{8'd76, 8'd21}: color_data = 12'hfc5;
			{8'd76, 8'd22}: color_data = 12'hfc5;
			{8'd76, 8'd23}: color_data = 12'hfc5;
			{8'd76, 8'd24}: color_data = 12'hfc5;
			{8'd76, 8'd25}: color_data = 12'hfc5;
			{8'd76, 8'd26}: color_data = 12'hfc5;
			{8'd76, 8'd27}: color_data = 12'hff7;
			{8'd76, 8'd56}: color_data = 12'h000;
			{8'd76, 8'd57}: color_data = 12'h601;
			{8'd76, 8'd58}: color_data = 12'hc11;
			{8'd76, 8'd59}: color_data = 12'hf12;
			{8'd76, 8'd60}: color_data = 12'he12;
			{8'd76, 8'd61}: color_data = 12'he12;
			{8'd76, 8'd62}: color_data = 12'he12;
			{8'd76, 8'd63}: color_data = 12'he12;
			{8'd76, 8'd64}: color_data = 12'he12;
			{8'd76, 8'd65}: color_data = 12'he12;
			{8'd76, 8'd66}: color_data = 12'hf12;
			{8'd76, 8'd67}: color_data = 12'hb11;
			{8'd76, 8'd68}: color_data = 12'h000;
			{8'd76, 8'd80}: color_data = 12'h777;
			{8'd76, 8'd81}: color_data = 12'hfff;
			{8'd76, 8'd82}: color_data = 12'hfff;
			{8'd76, 8'd83}: color_data = 12'hfff;
			{8'd76, 8'd84}: color_data = 12'hccc;
			{8'd76, 8'd85}: color_data = 12'heee;
			{8'd76, 8'd86}: color_data = 12'hfff;
			{8'd76, 8'd87}: color_data = 12'hccc;
			{8'd76, 8'd88}: color_data = 12'hbbb;
			{8'd76, 8'd89}: color_data = 12'hfff;
			{8'd76, 8'd90}: color_data = 12'h999;
			{8'd76, 8'd91}: color_data = 12'hfff;
			{8'd76, 8'd92}: color_data = 12'hfff;
			{8'd76, 8'd93}: color_data = 12'h778;
			{8'd76, 8'd94}: color_data = 12'h037;
			{8'd76, 8'd95}: color_data = 12'h047;
			{8'd76, 8'd96}: color_data = 12'h047;
			{8'd76, 8'd97}: color_data = 12'h047;
			{8'd76, 8'd98}: color_data = 12'h047;
			{8'd76, 8'd99}: color_data = 12'h05a;
			{8'd76, 8'd100}: color_data = 12'h06b;
			{8'd76, 8'd101}: color_data = 12'h06b;
			{8'd76, 8'd102}: color_data = 12'h06b;
			{8'd76, 8'd103}: color_data = 12'h06b;
			{8'd76, 8'd104}: color_data = 12'h06b;
			{8'd76, 8'd105}: color_data = 12'h06b;
			{8'd76, 8'd106}: color_data = 12'h06b;
			{8'd76, 8'd107}: color_data = 12'h06b;
			{8'd76, 8'd108}: color_data = 12'h06b;
			{8'd76, 8'd109}: color_data = 12'h06b;
			{8'd76, 8'd110}: color_data = 12'h06b;
			{8'd76, 8'd111}: color_data = 12'h06b;
			{8'd76, 8'd112}: color_data = 12'h06b;
			{8'd76, 8'd113}: color_data = 12'h06b;
			{8'd76, 8'd114}: color_data = 12'h06b;
			{8'd76, 8'd115}: color_data = 12'h06b;
			{8'd76, 8'd116}: color_data = 12'h06b;
			{8'd76, 8'd117}: color_data = 12'h06b;
			{8'd76, 8'd118}: color_data = 12'h06b;
			{8'd76, 8'd119}: color_data = 12'h047;
			{8'd76, 8'd120}: color_data = 12'h000;
			{8'd77, 8'd8}: color_data = 12'hfc4;
			{8'd77, 8'd9}: color_data = 12'hfc5;
			{8'd77, 8'd10}: color_data = 12'hfc5;
			{8'd77, 8'd11}: color_data = 12'hfc4;
			{8'd77, 8'd12}: color_data = 12'hea0;
			{8'd77, 8'd13}: color_data = 12'hea2;
			{8'd77, 8'd14}: color_data = 12'heb3;
			{8'd77, 8'd15}: color_data = 12'hfb4;
			{8'd77, 8'd16}: color_data = 12'hfc5;
			{8'd77, 8'd17}: color_data = 12'hfc5;
			{8'd77, 8'd18}: color_data = 12'hfc6;
			{8'd77, 8'd19}: color_data = 12'hfc6;
			{8'd77, 8'd20}: color_data = 12'hfc5;
			{8'd77, 8'd21}: color_data = 12'hfc5;
			{8'd77, 8'd22}: color_data = 12'hfc5;
			{8'd77, 8'd23}: color_data = 12'hfc5;
			{8'd77, 8'd24}: color_data = 12'hfc4;
			{8'd77, 8'd55}: color_data = 12'h000;
			{8'd77, 8'd56}: color_data = 12'h701;
			{8'd77, 8'd57}: color_data = 12'hd12;
			{8'd77, 8'd58}: color_data = 12'hf12;
			{8'd77, 8'd59}: color_data = 12'he12;
			{8'd77, 8'd60}: color_data = 12'he12;
			{8'd77, 8'd61}: color_data = 12'he12;
			{8'd77, 8'd62}: color_data = 12'he12;
			{8'd77, 8'd63}: color_data = 12'he12;
			{8'd77, 8'd64}: color_data = 12'he12;
			{8'd77, 8'd65}: color_data = 12'he12;
			{8'd77, 8'd66}: color_data = 12'hf12;
			{8'd77, 8'd67}: color_data = 12'h711;
			{8'd77, 8'd68}: color_data = 12'h211;
			{8'd77, 8'd69}: color_data = 12'h421;
			{8'd77, 8'd70}: color_data = 12'h421;
			{8'd77, 8'd71}: color_data = 12'h311;
			{8'd77, 8'd72}: color_data = 12'h100;
			{8'd77, 8'd73}: color_data = 12'h000;
			{8'd77, 8'd80}: color_data = 12'h666;
			{8'd77, 8'd81}: color_data = 12'hfff;
			{8'd77, 8'd82}: color_data = 12'hfff;
			{8'd77, 8'd83}: color_data = 12'hfff;
			{8'd77, 8'd84}: color_data = 12'heee;
			{8'd77, 8'd85}: color_data = 12'haaa;
			{8'd77, 8'd86}: color_data = 12'hfff;
			{8'd77, 8'd87}: color_data = 12'hfff;
			{8'd77, 8'd88}: color_data = 12'haaa;
			{8'd77, 8'd89}: color_data = 12'hbbb;
			{8'd77, 8'd90}: color_data = 12'hddd;
			{8'd77, 8'd91}: color_data = 12'h467;
			{8'd77, 8'd92}: color_data = 12'h358;
			{8'd77, 8'd93}: color_data = 12'h135;
			{8'd77, 8'd94}: color_data = 12'h256;
			{8'd77, 8'd95}: color_data = 12'h156;
			{8'd77, 8'd96}: color_data = 12'h05a;
			{8'd77, 8'd97}: color_data = 12'h06b;
			{8'd77, 8'd98}: color_data = 12'h05a;
			{8'd77, 8'd99}: color_data = 12'h036;
			{8'd77, 8'd100}: color_data = 12'h06b;
			{8'd77, 8'd101}: color_data = 12'h06b;
			{8'd77, 8'd102}: color_data = 12'h06b;
			{8'd77, 8'd103}: color_data = 12'h06b;
			{8'd77, 8'd104}: color_data = 12'h06b;
			{8'd77, 8'd105}: color_data = 12'h06b;
			{8'd77, 8'd106}: color_data = 12'h06b;
			{8'd77, 8'd107}: color_data = 12'h06b;
			{8'd77, 8'd108}: color_data = 12'h06b;
			{8'd77, 8'd109}: color_data = 12'h06b;
			{8'd77, 8'd110}: color_data = 12'h06b;
			{8'd77, 8'd111}: color_data = 12'h06b;
			{8'd77, 8'd112}: color_data = 12'h06b;
			{8'd77, 8'd113}: color_data = 12'h06b;
			{8'd77, 8'd114}: color_data = 12'h06b;
			{8'd77, 8'd115}: color_data = 12'h06b;
			{8'd77, 8'd116}: color_data = 12'h06b;
			{8'd77, 8'd117}: color_data = 12'h06b;
			{8'd77, 8'd118}: color_data = 12'h06b;
			{8'd77, 8'd119}: color_data = 12'h048;
			{8'd77, 8'd120}: color_data = 12'h000;
			{8'd78, 8'd8}: color_data = 12'hfc4;
			{8'd78, 8'd9}: color_data = 12'hfc5;
			{8'd78, 8'd10}: color_data = 12'hfc5;
			{8'd78, 8'd11}: color_data = 12'hfc4;
			{8'd78, 8'd12}: color_data = 12'hfc4;
			{8'd78, 8'd13}: color_data = 12'hfc4;
			{8'd78, 8'd14}: color_data = 12'hfc4;
			{8'd78, 8'd15}: color_data = 12'hfc5;
			{8'd78, 8'd16}: color_data = 12'hfc6;
			{8'd78, 8'd17}: color_data = 12'hfc5;
			{8'd78, 8'd18}: color_data = 12'hfc6;
			{8'd78, 8'd19}: color_data = 12'hfd7;
			{8'd78, 8'd20}: color_data = 12'hfd7;
			{8'd78, 8'd21}: color_data = 12'hfc5;
			{8'd78, 8'd54}: color_data = 12'h000;
			{8'd78, 8'd55}: color_data = 12'h701;
			{8'd78, 8'd56}: color_data = 12'hf12;
			{8'd78, 8'd57}: color_data = 12'hf12;
			{8'd78, 8'd58}: color_data = 12'he12;
			{8'd78, 8'd59}: color_data = 12'he12;
			{8'd78, 8'd60}: color_data = 12'he12;
			{8'd78, 8'd61}: color_data = 12'he12;
			{8'd78, 8'd62}: color_data = 12'he12;
			{8'd78, 8'd63}: color_data = 12'he12;
			{8'd78, 8'd64}: color_data = 12'he12;
			{8'd78, 8'd65}: color_data = 12'hf12;
			{8'd78, 8'd66}: color_data = 12'hc11;
			{8'd78, 8'd67}: color_data = 12'h631;
			{8'd78, 8'd68}: color_data = 12'h843;
			{8'd78, 8'd69}: color_data = 12'h843;
			{8'd78, 8'd70}: color_data = 12'h843;
			{8'd78, 8'd71}: color_data = 12'h843;
			{8'd78, 8'd72}: color_data = 12'h742;
			{8'd78, 8'd73}: color_data = 12'h321;
			{8'd78, 8'd74}: color_data = 12'h000;
			{8'd78, 8'd80}: color_data = 12'h222;
			{8'd78, 8'd81}: color_data = 12'hddd;
			{8'd78, 8'd82}: color_data = 12'hfff;
			{8'd78, 8'd83}: color_data = 12'hfff;
			{8'd78, 8'd84}: color_data = 12'hfff;
			{8'd78, 8'd85}: color_data = 12'hbbb;
			{8'd78, 8'd86}: color_data = 12'hbbb;
			{8'd78, 8'd87}: color_data = 12'hfff;
			{8'd78, 8'd88}: color_data = 12'hfff;
			{8'd78, 8'd89}: color_data = 12'hccc;
			{8'd78, 8'd90}: color_data = 12'h667;
			{8'd78, 8'd91}: color_data = 12'h036;
			{8'd78, 8'd92}: color_data = 12'h672;
			{8'd78, 8'd93}: color_data = 12'hdc0;
			{8'd78, 8'd94}: color_data = 12'hfe0;
			{8'd78, 8'd95}: color_data = 12'hfe0;
			{8'd78, 8'd96}: color_data = 12'h672;
			{8'd78, 8'd97}: color_data = 12'h05a;
			{8'd78, 8'd98}: color_data = 12'h06b;
			{8'd78, 8'd99}: color_data = 12'h047;
			{8'd78, 8'd100}: color_data = 12'h06a;
			{8'd78, 8'd101}: color_data = 12'h06b;
			{8'd78, 8'd102}: color_data = 12'h06b;
			{8'd78, 8'd103}: color_data = 12'h06b;
			{8'd78, 8'd104}: color_data = 12'h06b;
			{8'd78, 8'd105}: color_data = 12'h06b;
			{8'd78, 8'd106}: color_data = 12'h06b;
			{8'd78, 8'd107}: color_data = 12'h06b;
			{8'd78, 8'd108}: color_data = 12'h06b;
			{8'd78, 8'd109}: color_data = 12'h06b;
			{8'd78, 8'd110}: color_data = 12'h06b;
			{8'd78, 8'd111}: color_data = 12'h06b;
			{8'd78, 8'd112}: color_data = 12'h06b;
			{8'd78, 8'd113}: color_data = 12'h06b;
			{8'd78, 8'd114}: color_data = 12'h06b;
			{8'd78, 8'd115}: color_data = 12'h06b;
			{8'd78, 8'd116}: color_data = 12'h06b;
			{8'd78, 8'd117}: color_data = 12'h06b;
			{8'd78, 8'd118}: color_data = 12'h06b;
			{8'd78, 8'd119}: color_data = 12'h06a;
			{8'd78, 8'd120}: color_data = 12'h024;
			{8'd79, 8'd7}: color_data = 12'hfa5;
			{8'd79, 8'd8}: color_data = 12'hfc4;
			{8'd79, 8'd9}: color_data = 12'hfc5;
			{8'd79, 8'd10}: color_data = 12'hea1;
			{8'd79, 8'd11}: color_data = 12'hd90;
			{8'd79, 8'd12}: color_data = 12'hea0;
			{8'd79, 8'd13}: color_data = 12'hda0;
			{8'd79, 8'd14}: color_data = 12'hd90;
			{8'd79, 8'd15}: color_data = 12'hea0;
			{8'd79, 8'd16}: color_data = 12'hea2;
			{8'd79, 8'd17}: color_data = 12'heb3;
			{8'd79, 8'd18}: color_data = 12'hfc4;
			{8'd79, 8'd19}: color_data = 12'hfc5;
			{8'd79, 8'd20}: color_data = 12'hfc5;
			{8'd79, 8'd21}: color_data = 12'hfc4;
			{8'd79, 8'd22}: color_data = 12'hfc5;
			{8'd79, 8'd23}: color_data = 12'hfc5;
			{8'd79, 8'd24}: color_data = 12'hfc6;
			{8'd79, 8'd53}: color_data = 12'h000;
			{8'd79, 8'd54}: color_data = 12'h600;
			{8'd79, 8'd55}: color_data = 12'he12;
			{8'd79, 8'd56}: color_data = 12'he12;
			{8'd79, 8'd57}: color_data = 12'he12;
			{8'd79, 8'd58}: color_data = 12'he12;
			{8'd79, 8'd59}: color_data = 12'he12;
			{8'd79, 8'd60}: color_data = 12'he12;
			{8'd79, 8'd61}: color_data = 12'he12;
			{8'd79, 8'd62}: color_data = 12'he12;
			{8'd79, 8'd63}: color_data = 12'he12;
			{8'd79, 8'd64}: color_data = 12'he12;
			{8'd79, 8'd65}: color_data = 12'he12;
			{8'd79, 8'd66}: color_data = 12'h711;
			{8'd79, 8'd67}: color_data = 12'h842;
			{8'd79, 8'd68}: color_data = 12'h843;
			{8'd79, 8'd69}: color_data = 12'h842;
			{8'd79, 8'd70}: color_data = 12'h842;
			{8'd79, 8'd71}: color_data = 12'h842;
			{8'd79, 8'd72}: color_data = 12'h842;
			{8'd79, 8'd73}: color_data = 12'h843;
			{8'd79, 8'd74}: color_data = 12'h521;
			{8'd79, 8'd75}: color_data = 12'h000;
			{8'd79, 8'd78}: color_data = 12'h000;
			{8'd79, 8'd79}: color_data = 12'h000;
			{8'd79, 8'd80}: color_data = 12'h000;
			{8'd79, 8'd81}: color_data = 12'h755;
			{8'd79, 8'd82}: color_data = 12'heff;
			{8'd79, 8'd83}: color_data = 12'hfff;
			{8'd79, 8'd84}: color_data = 12'hfff;
			{8'd79, 8'd85}: color_data = 12'hfff;
			{8'd79, 8'd86}: color_data = 12'hbbb;
			{8'd79, 8'd87}: color_data = 12'haaa;
			{8'd79, 8'd88}: color_data = 12'hccc;
			{8'd79, 8'd89}: color_data = 12'h789;
			{8'd79, 8'd90}: color_data = 12'h047;
			{8'd79, 8'd91}: color_data = 12'h881;
			{8'd79, 8'd92}: color_data = 12'hff0;
			{8'd79, 8'd93}: color_data = 12'hff0;
			{8'd79, 8'd94}: color_data = 12'hff0;
			{8'd79, 8'd95}: color_data = 12'hff0;
			{8'd79, 8'd96}: color_data = 12'h891;
			{8'd79, 8'd97}: color_data = 12'h05a;
			{8'd79, 8'd98}: color_data = 12'h06b;
			{8'd79, 8'd99}: color_data = 12'h036;
			{8'd79, 8'd100}: color_data = 12'h06b;
			{8'd79, 8'd101}: color_data = 12'h06b;
			{8'd79, 8'd102}: color_data = 12'h06b;
			{8'd79, 8'd103}: color_data = 12'h06b;
			{8'd79, 8'd104}: color_data = 12'h06b;
			{8'd79, 8'd105}: color_data = 12'h06b;
			{8'd79, 8'd106}: color_data = 12'h06b;
			{8'd79, 8'd107}: color_data = 12'h06b;
			{8'd79, 8'd108}: color_data = 12'h06b;
			{8'd79, 8'd109}: color_data = 12'h06b;
			{8'd79, 8'd110}: color_data = 12'h06b;
			{8'd79, 8'd111}: color_data = 12'h06b;
			{8'd79, 8'd112}: color_data = 12'h06b;
			{8'd79, 8'd113}: color_data = 12'h06b;
			{8'd79, 8'd114}: color_data = 12'h06b;
			{8'd79, 8'd115}: color_data = 12'h06b;
			{8'd79, 8'd116}: color_data = 12'h06b;
			{8'd79, 8'd117}: color_data = 12'h06b;
			{8'd79, 8'd118}: color_data = 12'h06b;
			{8'd79, 8'd119}: color_data = 12'h06b;
			{8'd79, 8'd120}: color_data = 12'h048;
			{8'd79, 8'd121}: color_data = 12'h000;
			{8'd80, 8'd7}: color_data = 12'hfc6;
			{8'd80, 8'd8}: color_data = 12'hfc5;
			{8'd80, 8'd9}: color_data = 12'hfc5;
			{8'd80, 8'd10}: color_data = 12'hda0;
			{8'd80, 8'd11}: color_data = 12'hd90;
			{8'd80, 8'd12}: color_data = 12'hd90;
			{8'd80, 8'd13}: color_data = 12'hd90;
			{8'd80, 8'd14}: color_data = 12'hd90;
			{8'd80, 8'd15}: color_data = 12'hd90;
			{8'd80, 8'd16}: color_data = 12'hd90;
			{8'd80, 8'd17}: color_data = 12'hd90;
			{8'd80, 8'd18}: color_data = 12'hda0;
			{8'd80, 8'd19}: color_data = 12'hea1;
			{8'd80, 8'd20}: color_data = 12'hfb3;
			{8'd80, 8'd21}: color_data = 12'hfc4;
			{8'd80, 8'd22}: color_data = 12'hfc5;
			{8'd80, 8'd23}: color_data = 12'hfc5;
			{8'd80, 8'd24}: color_data = 12'hfc5;
			{8'd80, 8'd25}: color_data = 12'hfc5;
			{8'd80, 8'd53}: color_data = 12'h100;
			{8'd80, 8'd54}: color_data = 12'h911;
			{8'd80, 8'd55}: color_data = 12'h911;
			{8'd80, 8'd56}: color_data = 12'ha11;
			{8'd80, 8'd57}: color_data = 12'he12;
			{8'd80, 8'd58}: color_data = 12'he12;
			{8'd80, 8'd59}: color_data = 12'he12;
			{8'd80, 8'd60}: color_data = 12'he12;
			{8'd80, 8'd61}: color_data = 12'he12;
			{8'd80, 8'd62}: color_data = 12'he12;
			{8'd80, 8'd63}: color_data = 12'he12;
			{8'd80, 8'd64}: color_data = 12'hf12;
			{8'd80, 8'd65}: color_data = 12'ha11;
			{8'd80, 8'd66}: color_data = 12'h632;
			{8'd80, 8'd67}: color_data = 12'h843;
			{8'd80, 8'd68}: color_data = 12'h732;
			{8'd80, 8'd69}: color_data = 12'h642;
			{8'd80, 8'd70}: color_data = 12'h753;
			{8'd80, 8'd71}: color_data = 12'h754;
			{8'd80, 8'd72}: color_data = 12'h643;
			{8'd80, 8'd73}: color_data = 12'h632;
			{8'd80, 8'd74}: color_data = 12'h842;
			{8'd80, 8'd75}: color_data = 12'h532;
			{8'd80, 8'd76}: color_data = 12'h000;
			{8'd80, 8'd77}: color_data = 12'h000;
			{8'd80, 8'd78}: color_data = 12'h531;
			{8'd80, 8'd79}: color_data = 12'h321;
			{8'd80, 8'd80}: color_data = 12'h300;
			{8'd80, 8'd81}: color_data = 12'h811;
			{8'd80, 8'd82}: color_data = 12'h765;
			{8'd80, 8'd83}: color_data = 12'hbbb;
			{8'd80, 8'd84}: color_data = 12'hfff;
			{8'd80, 8'd85}: color_data = 12'hfff;
			{8'd80, 8'd86}: color_data = 12'hfff;
			{8'd80, 8'd87}: color_data = 12'h899;
			{8'd80, 8'd88}: color_data = 12'h047;
			{8'd80, 8'd89}: color_data = 12'h05a;
			{8'd80, 8'd90}: color_data = 12'h059;
			{8'd80, 8'd91}: color_data = 12'hcb0;
			{8'd80, 8'd92}: color_data = 12'hff0;
			{8'd80, 8'd93}: color_data = 12'hff0;
			{8'd80, 8'd94}: color_data = 12'hfe0;
			{8'd80, 8'd95}: color_data = 12'haa0;
			{8'd80, 8'd96}: color_data = 12'h157;
			{8'd80, 8'd97}: color_data = 12'h05a;
			{8'd80, 8'd98}: color_data = 12'h036;
			{8'd80, 8'd99}: color_data = 12'h059;
			{8'd80, 8'd100}: color_data = 12'h06b;
			{8'd80, 8'd101}: color_data = 12'h06b;
			{8'd80, 8'd102}: color_data = 12'h06b;
			{8'd80, 8'd103}: color_data = 12'h06b;
			{8'd80, 8'd104}: color_data = 12'h06b;
			{8'd80, 8'd105}: color_data = 12'h06b;
			{8'd80, 8'd106}: color_data = 12'h06b;
			{8'd80, 8'd107}: color_data = 12'h06b;
			{8'd80, 8'd108}: color_data = 12'h06b;
			{8'd80, 8'd109}: color_data = 12'h06b;
			{8'd80, 8'd110}: color_data = 12'h06b;
			{8'd80, 8'd111}: color_data = 12'h06b;
			{8'd80, 8'd112}: color_data = 12'h06b;
			{8'd80, 8'd113}: color_data = 12'h06b;
			{8'd80, 8'd114}: color_data = 12'h06b;
			{8'd80, 8'd115}: color_data = 12'h06b;
			{8'd80, 8'd116}: color_data = 12'h06b;
			{8'd80, 8'd117}: color_data = 12'h06b;
			{8'd80, 8'd118}: color_data = 12'h06b;
			{8'd80, 8'd119}: color_data = 12'h06b;
			{8'd80, 8'd120}: color_data = 12'h06b;
			{8'd80, 8'd121}: color_data = 12'h035;
			{8'd80, 8'd122}: color_data = 12'h000;
			{8'd81, 8'd7}: color_data = 12'hfc5;
			{8'd81, 8'd8}: color_data = 12'hfc5;
			{8'd81, 8'd9}: color_data = 12'hfc4;
			{8'd81, 8'd10}: color_data = 12'hd90;
			{8'd81, 8'd11}: color_data = 12'hd90;
			{8'd81, 8'd12}: color_data = 12'hd90;
			{8'd81, 8'd13}: color_data = 12'hd90;
			{8'd81, 8'd14}: color_data = 12'hd90;
			{8'd81, 8'd15}: color_data = 12'hd90;
			{8'd81, 8'd16}: color_data = 12'hd90;
			{8'd81, 8'd17}: color_data = 12'hd90;
			{8'd81, 8'd18}: color_data = 12'hd90;
			{8'd81, 8'd19}: color_data = 12'hd90;
			{8'd81, 8'd20}: color_data = 12'hd90;
			{8'd81, 8'd21}: color_data = 12'hd90;
			{8'd81, 8'd22}: color_data = 12'hea1;
			{8'd81, 8'd23}: color_data = 12'hfb3;
			{8'd81, 8'd24}: color_data = 12'hfc5;
			{8'd81, 8'd25}: color_data = 12'hfc5;
			{8'd81, 8'd49}: color_data = 12'h000;
			{8'd81, 8'd50}: color_data = 12'h100;
			{8'd81, 8'd51}: color_data = 12'h400;
			{8'd81, 8'd52}: color_data = 12'h701;
			{8'd81, 8'd53}: color_data = 12'ha11;
			{8'd81, 8'd54}: color_data = 12'hd12;
			{8'd81, 8'd55}: color_data = 12'he12;
			{8'd81, 8'd56}: color_data = 12'hf12;
			{8'd81, 8'd57}: color_data = 12'he12;
			{8'd81, 8'd58}: color_data = 12'he12;
			{8'd81, 8'd59}: color_data = 12'he12;
			{8'd81, 8'd60}: color_data = 12'he12;
			{8'd81, 8'd61}: color_data = 12'he12;
			{8'd81, 8'd62}: color_data = 12'he12;
			{8'd81, 8'd63}: color_data = 12'hf12;
			{8'd81, 8'd64}: color_data = 12'hd12;
			{8'd81, 8'd65}: color_data = 12'h621;
			{8'd81, 8'd66}: color_data = 12'h843;
			{8'd81, 8'd67}: color_data = 12'h632;
			{8'd81, 8'd68}: color_data = 12'h976;
			{8'd81, 8'd69}: color_data = 12'heca;
			{8'd81, 8'd70}: color_data = 12'hfdb;
			{8'd81, 8'd71}: color_data = 12'hfdb;
			{8'd81, 8'd72}: color_data = 12'heca;
			{8'd81, 8'd73}: color_data = 12'hb98;
			{8'd81, 8'd74}: color_data = 12'h754;
			{8'd81, 8'd75}: color_data = 12'h732;
			{8'd81, 8'd76}: color_data = 12'h521;
			{8'd81, 8'd77}: color_data = 12'h100;
			{8'd81, 8'd78}: color_data = 12'h842;
			{8'd81, 8'd79}: color_data = 12'h531;
			{8'd81, 8'd80}: color_data = 12'h100;
			{8'd81, 8'd81}: color_data = 12'h965;
			{8'd81, 8'd82}: color_data = 12'hc97;
			{8'd81, 8'd83}: color_data = 12'ha76;
			{8'd81, 8'd84}: color_data = 12'h876;
			{8'd81, 8'd85}: color_data = 12'h988;
			{8'd81, 8'd86}: color_data = 12'h899;
			{8'd81, 8'd87}: color_data = 12'h258;
			{8'd81, 8'd88}: color_data = 12'h06b;
			{8'd81, 8'd89}: color_data = 12'h06b;
			{8'd81, 8'd90}: color_data = 12'h06b;
			{8'd81, 8'd91}: color_data = 12'h256;
			{8'd81, 8'd92}: color_data = 12'h782;
			{8'd81, 8'd93}: color_data = 12'h782;
			{8'd81, 8'd94}: color_data = 12'h364;
			{8'd81, 8'd95}: color_data = 12'h048;
			{8'd81, 8'd96}: color_data = 12'h048;
			{8'd81, 8'd97}: color_data = 12'h047;
			{8'd81, 8'd98}: color_data = 12'h05a;
			{8'd81, 8'd99}: color_data = 12'h06b;
			{8'd81, 8'd100}: color_data = 12'h06b;
			{8'd81, 8'd101}: color_data = 12'h06b;
			{8'd81, 8'd102}: color_data = 12'h06b;
			{8'd81, 8'd103}: color_data = 12'h06b;
			{8'd81, 8'd104}: color_data = 12'h06b;
			{8'd81, 8'd105}: color_data = 12'h06b;
			{8'd81, 8'd106}: color_data = 12'h06b;
			{8'd81, 8'd107}: color_data = 12'h06b;
			{8'd81, 8'd108}: color_data = 12'h06b;
			{8'd81, 8'd109}: color_data = 12'h06b;
			{8'd81, 8'd110}: color_data = 12'h06b;
			{8'd81, 8'd111}: color_data = 12'h06b;
			{8'd81, 8'd112}: color_data = 12'h06b;
			{8'd81, 8'd113}: color_data = 12'h06b;
			{8'd81, 8'd114}: color_data = 12'h06b;
			{8'd81, 8'd115}: color_data = 12'h06b;
			{8'd81, 8'd116}: color_data = 12'h06b;
			{8'd81, 8'd117}: color_data = 12'h06b;
			{8'd81, 8'd118}: color_data = 12'h06b;
			{8'd81, 8'd119}: color_data = 12'h06b;
			{8'd81, 8'd120}: color_data = 12'h06b;
			{8'd81, 8'd121}: color_data = 12'h058;
			{8'd81, 8'd122}: color_data = 12'h000;
			{8'd82, 8'd7}: color_data = 12'hfc5;
			{8'd82, 8'd8}: color_data = 12'hfc5;
			{8'd82, 8'd9}: color_data = 12'heb3;
			{8'd82, 8'd10}: color_data = 12'hd90;
			{8'd82, 8'd11}: color_data = 12'hd90;
			{8'd82, 8'd12}: color_data = 12'hd90;
			{8'd82, 8'd13}: color_data = 12'hd90;
			{8'd82, 8'd14}: color_data = 12'hd90;
			{8'd82, 8'd15}: color_data = 12'hd90;
			{8'd82, 8'd16}: color_data = 12'hd90;
			{8'd82, 8'd17}: color_data = 12'hd90;
			{8'd82, 8'd18}: color_data = 12'hd90;
			{8'd82, 8'd19}: color_data = 12'hd90;
			{8'd82, 8'd20}: color_data = 12'hd90;
			{8'd82, 8'd21}: color_data = 12'hd90;
			{8'd82, 8'd22}: color_data = 12'hd90;
			{8'd82, 8'd23}: color_data = 12'hea1;
			{8'd82, 8'd24}: color_data = 12'hfc5;
			{8'd82, 8'd25}: color_data = 12'hfc5;
			{8'd82, 8'd46}: color_data = 12'h000;
			{8'd82, 8'd47}: color_data = 12'h100;
			{8'd82, 8'd48}: color_data = 12'h500;
			{8'd82, 8'd49}: color_data = 12'h911;
			{8'd82, 8'd50}: color_data = 12'hc11;
			{8'd82, 8'd51}: color_data = 12'he12;
			{8'd82, 8'd52}: color_data = 12'hf12;
			{8'd82, 8'd53}: color_data = 12'hf12;
			{8'd82, 8'd54}: color_data = 12'hf12;
			{8'd82, 8'd55}: color_data = 12'he12;
			{8'd82, 8'd56}: color_data = 12'he12;
			{8'd82, 8'd57}: color_data = 12'he12;
			{8'd82, 8'd58}: color_data = 12'he12;
			{8'd82, 8'd59}: color_data = 12'he12;
			{8'd82, 8'd60}: color_data = 12'he12;
			{8'd82, 8'd61}: color_data = 12'he12;
			{8'd82, 8'd62}: color_data = 12'he12;
			{8'd82, 8'd63}: color_data = 12'hf12;
			{8'd82, 8'd64}: color_data = 12'h811;
			{8'd82, 8'd65}: color_data = 12'h742;
			{8'd82, 8'd66}: color_data = 12'h742;
			{8'd82, 8'd67}: color_data = 12'h865;
			{8'd82, 8'd68}: color_data = 12'hfdb;
			{8'd82, 8'd69}: color_data = 12'hfdb;
			{8'd82, 8'd70}: color_data = 12'hfdb;
			{8'd82, 8'd71}: color_data = 12'hfda;
			{8'd82, 8'd72}: color_data = 12'hfdb;
			{8'd82, 8'd73}: color_data = 12'hfdb;
			{8'd82, 8'd74}: color_data = 12'hfdb;
			{8'd82, 8'd75}: color_data = 12'ha87;
			{8'd82, 8'd76}: color_data = 12'h632;
			{8'd82, 8'd77}: color_data = 12'h531;
			{8'd82, 8'd78}: color_data = 12'h843;
			{8'd82, 8'd79}: color_data = 12'h632;
			{8'd82, 8'd80}: color_data = 12'h421;
			{8'd82, 8'd81}: color_data = 12'hb87;
			{8'd82, 8'd82}: color_data = 12'hc97;
			{8'd82, 8'd83}: color_data = 12'hd97;
			{8'd82, 8'd84}: color_data = 12'h975;
			{8'd82, 8'd85}: color_data = 12'h036;
			{8'd82, 8'd86}: color_data = 12'h05a;
			{8'd82, 8'd87}: color_data = 12'h06b;
			{8'd82, 8'd88}: color_data = 12'h06b;
			{8'd82, 8'd89}: color_data = 12'h06b;
			{8'd82, 8'd90}: color_data = 12'h06b;
			{8'd82, 8'd91}: color_data = 12'h06b;
			{8'd82, 8'd92}: color_data = 12'h05b;
			{8'd82, 8'd93}: color_data = 12'h049;
			{8'd82, 8'd94}: color_data = 12'h037;
			{8'd82, 8'd95}: color_data = 12'h047;
			{8'd82, 8'd96}: color_data = 12'h059;
			{8'd82, 8'd97}: color_data = 12'h06b;
			{8'd82, 8'd98}: color_data = 12'h06b;
			{8'd82, 8'd99}: color_data = 12'h06b;
			{8'd82, 8'd100}: color_data = 12'h06b;
			{8'd82, 8'd101}: color_data = 12'h06b;
			{8'd82, 8'd102}: color_data = 12'h06b;
			{8'd82, 8'd103}: color_data = 12'h06b;
			{8'd82, 8'd104}: color_data = 12'h06b;
			{8'd82, 8'd105}: color_data = 12'h06b;
			{8'd82, 8'd106}: color_data = 12'h06b;
			{8'd82, 8'd107}: color_data = 12'h06b;
			{8'd82, 8'd108}: color_data = 12'h06b;
			{8'd82, 8'd109}: color_data = 12'h06b;
			{8'd82, 8'd110}: color_data = 12'h06b;
			{8'd82, 8'd111}: color_data = 12'h06b;
			{8'd82, 8'd112}: color_data = 12'h06b;
			{8'd82, 8'd113}: color_data = 12'h06b;
			{8'd82, 8'd114}: color_data = 12'h06b;
			{8'd82, 8'd115}: color_data = 12'h06b;
			{8'd82, 8'd116}: color_data = 12'h06b;
			{8'd82, 8'd117}: color_data = 12'h06b;
			{8'd82, 8'd118}: color_data = 12'h06b;
			{8'd82, 8'd119}: color_data = 12'h06b;
			{8'd82, 8'd120}: color_data = 12'h06b;
			{8'd82, 8'd121}: color_data = 12'h06b;
			{8'd82, 8'd122}: color_data = 12'h024;
			{8'd83, 8'd7}: color_data = 12'hfc5;
			{8'd83, 8'd8}: color_data = 12'hfc5;
			{8'd83, 8'd9}: color_data = 12'heb2;
			{8'd83, 8'd10}: color_data = 12'hd90;
			{8'd83, 8'd11}: color_data = 12'hd90;
			{8'd83, 8'd12}: color_data = 12'hd90;
			{8'd83, 8'd13}: color_data = 12'hd90;
			{8'd83, 8'd14}: color_data = 12'hea1;
			{8'd83, 8'd15}: color_data = 12'hd90;
			{8'd83, 8'd16}: color_data = 12'hd90;
			{8'd83, 8'd17}: color_data = 12'hd90;
			{8'd83, 8'd18}: color_data = 12'hd90;
			{8'd83, 8'd19}: color_data = 12'hd90;
			{8'd83, 8'd20}: color_data = 12'hd90;
			{8'd83, 8'd21}: color_data = 12'hd90;
			{8'd83, 8'd22}: color_data = 12'hd90;
			{8'd83, 8'd23}: color_data = 12'heb2;
			{8'd83, 8'd24}: color_data = 12'hfc6;
			{8'd83, 8'd25}: color_data = 12'hfc5;
			{8'd83, 8'd44}: color_data = 12'h000;
			{8'd83, 8'd45}: color_data = 12'h300;
			{8'd83, 8'd46}: color_data = 12'h701;
			{8'd83, 8'd47}: color_data = 12'hb11;
			{8'd83, 8'd48}: color_data = 12'he12;
			{8'd83, 8'd49}: color_data = 12'hf12;
			{8'd83, 8'd50}: color_data = 12'hf12;
			{8'd83, 8'd51}: color_data = 12'he12;
			{8'd83, 8'd52}: color_data = 12'he12;
			{8'd83, 8'd53}: color_data = 12'he12;
			{8'd83, 8'd54}: color_data = 12'he12;
			{8'd83, 8'd55}: color_data = 12'he12;
			{8'd83, 8'd56}: color_data = 12'he12;
			{8'd83, 8'd57}: color_data = 12'he12;
			{8'd83, 8'd58}: color_data = 12'he12;
			{8'd83, 8'd59}: color_data = 12'he12;
			{8'd83, 8'd60}: color_data = 12'he12;
			{8'd83, 8'd61}: color_data = 12'he12;
			{8'd83, 8'd62}: color_data = 12'hf12;
			{8'd83, 8'd63}: color_data = 12'hb11;
			{8'd83, 8'd64}: color_data = 12'h632;
			{8'd83, 8'd65}: color_data = 12'h843;
			{8'd83, 8'd66}: color_data = 12'h732;
			{8'd83, 8'd67}: color_data = 12'ha87;
			{8'd83, 8'd68}: color_data = 12'hfdb;
			{8'd83, 8'd69}: color_data = 12'hfca;
			{8'd83, 8'd70}: color_data = 12'hfca;
			{8'd83, 8'd71}: color_data = 12'hfdb;
			{8'd83, 8'd72}: color_data = 12'hfdb;
			{8'd83, 8'd73}: color_data = 12'hfda;
			{8'd83, 8'd74}: color_data = 12'hfdb;
			{8'd83, 8'd75}: color_data = 12'hfdb;
			{8'd83, 8'd76}: color_data = 12'hda9;
			{8'd83, 8'd77}: color_data = 12'h643;
			{8'd83, 8'd78}: color_data = 12'h842;
			{8'd83, 8'd79}: color_data = 12'h843;
			{8'd83, 8'd80}: color_data = 12'h632;
			{8'd83, 8'd81}: color_data = 12'ha76;
			{8'd83, 8'd82}: color_data = 12'hd97;
			{8'd83, 8'd83}: color_data = 12'h975;
			{8'd83, 8'd84}: color_data = 12'h047;
			{8'd83, 8'd85}: color_data = 12'h06b;
			{8'd83, 8'd86}: color_data = 12'h06b;
			{8'd83, 8'd87}: color_data = 12'h06b;
			{8'd83, 8'd88}: color_data = 12'h06b;
			{8'd83, 8'd89}: color_data = 12'h06b;
			{8'd83, 8'd90}: color_data = 12'h06b;
			{8'd83, 8'd91}: color_data = 12'h048;
			{8'd83, 8'd92}: color_data = 12'h125;
			{8'd83, 8'd93}: color_data = 12'h047;
			{8'd83, 8'd94}: color_data = 12'h05a;
			{8'd83, 8'd95}: color_data = 12'h06b;
			{8'd83, 8'd96}: color_data = 12'h06b;
			{8'd83, 8'd97}: color_data = 12'h06b;
			{8'd83, 8'd98}: color_data = 12'h06b;
			{8'd83, 8'd99}: color_data = 12'h06b;
			{8'd83, 8'd100}: color_data = 12'h06b;
			{8'd83, 8'd101}: color_data = 12'h06b;
			{8'd83, 8'd102}: color_data = 12'h06b;
			{8'd83, 8'd103}: color_data = 12'h06b;
			{8'd83, 8'd104}: color_data = 12'h06b;
			{8'd83, 8'd105}: color_data = 12'h06b;
			{8'd83, 8'd106}: color_data = 12'h06b;
			{8'd83, 8'd107}: color_data = 12'h06b;
			{8'd83, 8'd108}: color_data = 12'h06b;
			{8'd83, 8'd109}: color_data = 12'h06b;
			{8'd83, 8'd110}: color_data = 12'h06b;
			{8'd83, 8'd111}: color_data = 12'h06b;
			{8'd83, 8'd112}: color_data = 12'h06b;
			{8'd83, 8'd113}: color_data = 12'h06b;
			{8'd83, 8'd114}: color_data = 12'h06b;
			{8'd83, 8'd115}: color_data = 12'h06b;
			{8'd83, 8'd116}: color_data = 12'h06b;
			{8'd83, 8'd117}: color_data = 12'h06b;
			{8'd83, 8'd118}: color_data = 12'h06b;
			{8'd83, 8'd119}: color_data = 12'h06b;
			{8'd83, 8'd120}: color_data = 12'h06b;
			{8'd83, 8'd121}: color_data = 12'h06b;
			{8'd83, 8'd122}: color_data = 12'h037;
			{8'd83, 8'd123}: color_data = 12'h000;
			{8'd84, 8'd7}: color_data = 12'hfc5;
			{8'd84, 8'd8}: color_data = 12'hfc5;
			{8'd84, 8'd9}: color_data = 12'hea1;
			{8'd84, 8'd10}: color_data = 12'hd90;
			{8'd84, 8'd11}: color_data = 12'hd90;
			{8'd84, 8'd12}: color_data = 12'hd90;
			{8'd84, 8'd13}: color_data = 12'hea2;
			{8'd84, 8'd14}: color_data = 12'hfc4;
			{8'd84, 8'd15}: color_data = 12'hd90;
			{8'd84, 8'd16}: color_data = 12'hd90;
			{8'd84, 8'd17}: color_data = 12'hd90;
			{8'd84, 8'd18}: color_data = 12'hea0;
			{8'd84, 8'd19}: color_data = 12'hd90;
			{8'd84, 8'd20}: color_data = 12'hd90;
			{8'd84, 8'd21}: color_data = 12'hd90;
			{8'd84, 8'd22}: color_data = 12'hd90;
			{8'd84, 8'd23}: color_data = 12'hfb3;
			{8'd84, 8'd24}: color_data = 12'hfc5;
			{8'd84, 8'd25}: color_data = 12'hfc5;
			{8'd84, 8'd42}: color_data = 12'h000;
			{8'd84, 8'd43}: color_data = 12'h300;
			{8'd84, 8'd44}: color_data = 12'h811;
			{8'd84, 8'd45}: color_data = 12'hd12;
			{8'd84, 8'd46}: color_data = 12'hf12;
			{8'd84, 8'd47}: color_data = 12'hf12;
			{8'd84, 8'd48}: color_data = 12'he12;
			{8'd84, 8'd49}: color_data = 12'he12;
			{8'd84, 8'd50}: color_data = 12'he12;
			{8'd84, 8'd51}: color_data = 12'he12;
			{8'd84, 8'd52}: color_data = 12'he12;
			{8'd84, 8'd53}: color_data = 12'he12;
			{8'd84, 8'd54}: color_data = 12'he12;
			{8'd84, 8'd55}: color_data = 12'he12;
			{8'd84, 8'd56}: color_data = 12'he12;
			{8'd84, 8'd57}: color_data = 12'he12;
			{8'd84, 8'd58}: color_data = 12'he12;
			{8'd84, 8'd59}: color_data = 12'he12;
			{8'd84, 8'd60}: color_data = 12'he12;
			{8'd84, 8'd61}: color_data = 12'hf12;
			{8'd84, 8'd62}: color_data = 12'hd12;
			{8'd84, 8'd63}: color_data = 12'h621;
			{8'd84, 8'd64}: color_data = 12'h843;
			{8'd84, 8'd65}: color_data = 12'h842;
			{8'd84, 8'd66}: color_data = 12'h742;
			{8'd84, 8'd67}: color_data = 12'h976;
			{8'd84, 8'd68}: color_data = 12'hfdb;
			{8'd84, 8'd69}: color_data = 12'ha87;
			{8'd84, 8'd70}: color_data = 12'hdb9;
			{8'd84, 8'd71}: color_data = 12'hca8;
			{8'd84, 8'd72}: color_data = 12'hdb9;
			{8'd84, 8'd73}: color_data = 12'hfca;
			{8'd84, 8'd74}: color_data = 12'hfda;
			{8'd84, 8'd75}: color_data = 12'hfda;
			{8'd84, 8'd76}: color_data = 12'hfdb;
			{8'd84, 8'd77}: color_data = 12'hca8;
			{8'd84, 8'd78}: color_data = 12'h632;
			{8'd84, 8'd79}: color_data = 12'h843;
			{8'd84, 8'd80}: color_data = 12'h632;
			{8'd84, 8'd81}: color_data = 12'ha76;
			{8'd84, 8'd82}: color_data = 12'ha75;
			{8'd84, 8'd83}: color_data = 12'h147;
			{8'd84, 8'd84}: color_data = 12'h06b;
			{8'd84, 8'd85}: color_data = 12'h06b;
			{8'd84, 8'd86}: color_data = 12'h06b;
			{8'd84, 8'd87}: color_data = 12'h06b;
			{8'd84, 8'd88}: color_data = 12'h05a;
			{8'd84, 8'd89}: color_data = 12'h147;
			{8'd84, 8'd90}: color_data = 12'h623;
			{8'd84, 8'd91}: color_data = 12'hc11;
			{8'd84, 8'd92}: color_data = 12'h712;
			{8'd84, 8'd93}: color_data = 12'h06b;
			{8'd84, 8'd94}: color_data = 12'h06b;
			{8'd84, 8'd95}: color_data = 12'h06b;
			{8'd84, 8'd96}: color_data = 12'h06b;
			{8'd84, 8'd97}: color_data = 12'h06b;
			{8'd84, 8'd98}: color_data = 12'h06b;
			{8'd84, 8'd99}: color_data = 12'h06b;
			{8'd84, 8'd100}: color_data = 12'h06b;
			{8'd84, 8'd101}: color_data = 12'h06b;
			{8'd84, 8'd102}: color_data = 12'h06b;
			{8'd84, 8'd103}: color_data = 12'h06b;
			{8'd84, 8'd104}: color_data = 12'h06b;
			{8'd84, 8'd105}: color_data = 12'h06b;
			{8'd84, 8'd106}: color_data = 12'h06b;
			{8'd84, 8'd107}: color_data = 12'h06b;
			{8'd84, 8'd108}: color_data = 12'h06b;
			{8'd84, 8'd109}: color_data = 12'h06b;
			{8'd84, 8'd110}: color_data = 12'h06b;
			{8'd84, 8'd111}: color_data = 12'h06b;
			{8'd84, 8'd112}: color_data = 12'h06b;
			{8'd84, 8'd113}: color_data = 12'h06b;
			{8'd84, 8'd114}: color_data = 12'h06b;
			{8'd84, 8'd115}: color_data = 12'h06b;
			{8'd84, 8'd116}: color_data = 12'h06b;
			{8'd84, 8'd117}: color_data = 12'h06b;
			{8'd84, 8'd118}: color_data = 12'h06b;
			{8'd84, 8'd119}: color_data = 12'h06b;
			{8'd84, 8'd120}: color_data = 12'h06b;
			{8'd84, 8'd121}: color_data = 12'h06b;
			{8'd84, 8'd122}: color_data = 12'h059;
			{8'd84, 8'd123}: color_data = 12'h001;
			{8'd85, 8'd7}: color_data = 12'hfc4;
			{8'd85, 8'd8}: color_data = 12'hfc4;
			{8'd85, 8'd9}: color_data = 12'hd90;
			{8'd85, 8'd10}: color_data = 12'hd90;
			{8'd85, 8'd11}: color_data = 12'hd90;
			{8'd85, 8'd12}: color_data = 12'hd90;
			{8'd85, 8'd13}: color_data = 12'hfc4;
			{8'd85, 8'd14}: color_data = 12'hfc4;
			{8'd85, 8'd15}: color_data = 12'hd90;
			{8'd85, 8'd16}: color_data = 12'hd90;
			{8'd85, 8'd17}: color_data = 12'hd90;
			{8'd85, 8'd18}: color_data = 12'hfb3;
			{8'd85, 8'd19}: color_data = 12'hea1;
			{8'd85, 8'd20}: color_data = 12'hd90;
			{8'd85, 8'd21}: color_data = 12'hd90;
			{8'd85, 8'd22}: color_data = 12'hd90;
			{8'd85, 8'd23}: color_data = 12'hfc4;
			{8'd85, 8'd24}: color_data = 12'hfc5;
			{8'd85, 8'd25}: color_data = 12'hfc5;
			{8'd85, 8'd41}: color_data = 12'h000;
			{8'd85, 8'd42}: color_data = 12'h701;
			{8'd85, 8'd43}: color_data = 12'hd12;
			{8'd85, 8'd44}: color_data = 12'hf12;
			{8'd85, 8'd45}: color_data = 12'hf12;
			{8'd85, 8'd46}: color_data = 12'he12;
			{8'd85, 8'd47}: color_data = 12'he12;
			{8'd85, 8'd48}: color_data = 12'he12;
			{8'd85, 8'd49}: color_data = 12'he12;
			{8'd85, 8'd50}: color_data = 12'he12;
			{8'd85, 8'd51}: color_data = 12'he12;
			{8'd85, 8'd52}: color_data = 12'he12;
			{8'd85, 8'd53}: color_data = 12'he12;
			{8'd85, 8'd54}: color_data = 12'he12;
			{8'd85, 8'd55}: color_data = 12'he12;
			{8'd85, 8'd56}: color_data = 12'he12;
			{8'd85, 8'd57}: color_data = 12'he12;
			{8'd85, 8'd58}: color_data = 12'he12;
			{8'd85, 8'd59}: color_data = 12'he12;
			{8'd85, 8'd60}: color_data = 12'he12;
			{8'd85, 8'd61}: color_data = 12'hf12;
			{8'd85, 8'd62}: color_data = 12'h711;
			{8'd85, 8'd63}: color_data = 12'h742;
			{8'd85, 8'd64}: color_data = 12'h843;
			{8'd85, 8'd65}: color_data = 12'h842;
			{8'd85, 8'd66}: color_data = 12'h842;
			{8'd85, 8'd67}: color_data = 12'h754;
			{8'd85, 8'd68}: color_data = 12'hfca;
			{8'd85, 8'd69}: color_data = 12'h986;
			{8'd85, 8'd70}: color_data = 12'ha87;
			{8'd85, 8'd71}: color_data = 12'hb98;
			{8'd85, 8'd72}: color_data = 12'hb98;
			{8'd85, 8'd73}: color_data = 12'hfca;
			{8'd85, 8'd74}: color_data = 12'hfdb;
			{8'd85, 8'd75}: color_data = 12'hfda;
			{8'd85, 8'd76}: color_data = 12'hfdb;
			{8'd85, 8'd77}: color_data = 12'hfca;
			{8'd85, 8'd78}: color_data = 12'h743;
			{8'd85, 8'd79}: color_data = 12'h842;
			{8'd85, 8'd80}: color_data = 12'h642;
			{8'd85, 8'd81}: color_data = 12'h965;
			{8'd85, 8'd82}: color_data = 12'h147;
			{8'd85, 8'd83}: color_data = 12'h06b;
			{8'd85, 8'd84}: color_data = 12'h06b;
			{8'd85, 8'd85}: color_data = 12'h06b;
			{8'd85, 8'd86}: color_data = 12'h05a;
			{8'd85, 8'd87}: color_data = 12'h136;
			{8'd85, 8'd88}: color_data = 12'h712;
			{8'd85, 8'd89}: color_data = 12'hd11;
			{8'd85, 8'd90}: color_data = 12'hf12;
			{8'd85, 8'd91}: color_data = 12'hf12;
			{8'd85, 8'd92}: color_data = 12'h812;
			{8'd85, 8'd93}: color_data = 12'h06a;
			{8'd85, 8'd94}: color_data = 12'h06b;
			{8'd85, 8'd95}: color_data = 12'h06b;
			{8'd85, 8'd96}: color_data = 12'h06b;
			{8'd85, 8'd97}: color_data = 12'h06b;
			{8'd85, 8'd98}: color_data = 12'h06b;
			{8'd85, 8'd99}: color_data = 12'h06b;
			{8'd85, 8'd100}: color_data = 12'h06b;
			{8'd85, 8'd101}: color_data = 12'h06b;
			{8'd85, 8'd102}: color_data = 12'h06b;
			{8'd85, 8'd103}: color_data = 12'h06b;
			{8'd85, 8'd104}: color_data = 12'h06b;
			{8'd85, 8'd105}: color_data = 12'h06b;
			{8'd85, 8'd106}: color_data = 12'h06b;
			{8'd85, 8'd107}: color_data = 12'h06b;
			{8'd85, 8'd108}: color_data = 12'h06b;
			{8'd85, 8'd109}: color_data = 12'h06b;
			{8'd85, 8'd110}: color_data = 12'h06b;
			{8'd85, 8'd111}: color_data = 12'h06b;
			{8'd85, 8'd112}: color_data = 12'h06b;
			{8'd85, 8'd113}: color_data = 12'h06b;
			{8'd85, 8'd114}: color_data = 12'h06b;
			{8'd85, 8'd115}: color_data = 12'h06b;
			{8'd85, 8'd116}: color_data = 12'h06b;
			{8'd85, 8'd117}: color_data = 12'h06b;
			{8'd85, 8'd118}: color_data = 12'h06b;
			{8'd85, 8'd119}: color_data = 12'h06b;
			{8'd85, 8'd120}: color_data = 12'h06b;
			{8'd85, 8'd121}: color_data = 12'h06b;
			{8'd85, 8'd122}: color_data = 12'h06b;
			{8'd85, 8'd123}: color_data = 12'h013;
			{8'd85, 8'd124}: color_data = 12'h000;
			{8'd85, 8'd145}: color_data = 12'h000;
			{8'd85, 8'd146}: color_data = 12'h000;
			{8'd85, 8'd147}: color_data = 12'h000;
			{8'd86, 8'd7}: color_data = 12'hfc4;
			{8'd86, 8'd8}: color_data = 12'hfc4;
			{8'd86, 8'd9}: color_data = 12'hd90;
			{8'd86, 8'd10}: color_data = 12'hd90;
			{8'd86, 8'd11}: color_data = 12'hd90;
			{8'd86, 8'd12}: color_data = 12'hea0;
			{8'd86, 8'd13}: color_data = 12'hfc5;
			{8'd86, 8'd14}: color_data = 12'heb3;
			{8'd86, 8'd15}: color_data = 12'hd90;
			{8'd86, 8'd16}: color_data = 12'hd90;
			{8'd86, 8'd17}: color_data = 12'hea0;
			{8'd86, 8'd18}: color_data = 12'hfc5;
			{8'd86, 8'd19}: color_data = 12'hea1;
			{8'd86, 8'd20}: color_data = 12'hd90;
			{8'd86, 8'd21}: color_data = 12'hd90;
			{8'd86, 8'd22}: color_data = 12'hda0;
			{8'd86, 8'd23}: color_data = 12'hfc5;
			{8'd86, 8'd24}: color_data = 12'hfc5;
			{8'd86, 8'd25}: color_data = 12'hfc4;
			{8'd86, 8'd39}: color_data = 12'h000;
			{8'd86, 8'd40}: color_data = 12'h300;
			{8'd86, 8'd41}: color_data = 12'ha11;
			{8'd86, 8'd42}: color_data = 12'hf12;
			{8'd86, 8'd43}: color_data = 12'hf12;
			{8'd86, 8'd44}: color_data = 12'he12;
			{8'd86, 8'd45}: color_data = 12'he12;
			{8'd86, 8'd46}: color_data = 12'he12;
			{8'd86, 8'd47}: color_data = 12'he12;
			{8'd86, 8'd48}: color_data = 12'he12;
			{8'd86, 8'd49}: color_data = 12'he12;
			{8'd86, 8'd50}: color_data = 12'he12;
			{8'd86, 8'd51}: color_data = 12'he12;
			{8'd86, 8'd52}: color_data = 12'he12;
			{8'd86, 8'd53}: color_data = 12'he12;
			{8'd86, 8'd54}: color_data = 12'he12;
			{8'd86, 8'd55}: color_data = 12'he12;
			{8'd86, 8'd56}: color_data = 12'he12;
			{8'd86, 8'd57}: color_data = 12'he12;
			{8'd86, 8'd58}: color_data = 12'he12;
			{8'd86, 8'd59}: color_data = 12'he12;
			{8'd86, 8'd60}: color_data = 12'hf12;
			{8'd86, 8'd61}: color_data = 12'ha11;
			{8'd86, 8'd62}: color_data = 12'h632;
			{8'd86, 8'd63}: color_data = 12'h843;
			{8'd86, 8'd64}: color_data = 12'h842;
			{8'd86, 8'd65}: color_data = 12'h842;
			{8'd86, 8'd66}: color_data = 12'h842;
			{8'd86, 8'd67}: color_data = 12'h642;
			{8'd86, 8'd68}: color_data = 12'heb9;
			{8'd86, 8'd69}: color_data = 12'h765;
			{8'd86, 8'd70}: color_data = 12'hb98;
			{8'd86, 8'd71}: color_data = 12'hfdb;
			{8'd86, 8'd72}: color_data = 12'hfdb;
			{8'd86, 8'd73}: color_data = 12'hfdb;
			{8'd86, 8'd74}: color_data = 12'hfda;
			{8'd86, 8'd75}: color_data = 12'hfda;
			{8'd86, 8'd76}: color_data = 12'hfda;
			{8'd86, 8'd77}: color_data = 12'hfdb;
			{8'd86, 8'd78}: color_data = 12'h754;
			{8'd86, 8'd79}: color_data = 12'h632;
			{8'd86, 8'd80}: color_data = 12'h432;
			{8'd86, 8'd81}: color_data = 12'h147;
			{8'd86, 8'd82}: color_data = 12'h06b;
			{8'd86, 8'd83}: color_data = 12'h06b;
			{8'd86, 8'd84}: color_data = 12'h06a;
			{8'd86, 8'd85}: color_data = 12'h136;
			{8'd86, 8'd86}: color_data = 12'h812;
			{8'd86, 8'd87}: color_data = 12'hd11;
			{8'd86, 8'd88}: color_data = 12'hf12;
			{8'd86, 8'd89}: color_data = 12'hf12;
			{8'd86, 8'd90}: color_data = 12'he12;
			{8'd86, 8'd91}: color_data = 12'hf12;
			{8'd86, 8'd92}: color_data = 12'h812;
			{8'd86, 8'd93}: color_data = 12'h05a;
			{8'd86, 8'd94}: color_data = 12'h06b;
			{8'd86, 8'd95}: color_data = 12'h06b;
			{8'd86, 8'd96}: color_data = 12'h06b;
			{8'd86, 8'd97}: color_data = 12'h06b;
			{8'd86, 8'd98}: color_data = 12'h06b;
			{8'd86, 8'd99}: color_data = 12'h06b;
			{8'd86, 8'd100}: color_data = 12'h06b;
			{8'd86, 8'd101}: color_data = 12'h06b;
			{8'd86, 8'd102}: color_data = 12'h06b;
			{8'd86, 8'd103}: color_data = 12'h06b;
			{8'd86, 8'd104}: color_data = 12'h06b;
			{8'd86, 8'd105}: color_data = 12'h06b;
			{8'd86, 8'd106}: color_data = 12'h06b;
			{8'd86, 8'd107}: color_data = 12'h06b;
			{8'd86, 8'd108}: color_data = 12'h06b;
			{8'd86, 8'd109}: color_data = 12'h06b;
			{8'd86, 8'd110}: color_data = 12'h06b;
			{8'd86, 8'd111}: color_data = 12'h06b;
			{8'd86, 8'd112}: color_data = 12'h06b;
			{8'd86, 8'd113}: color_data = 12'h06b;
			{8'd86, 8'd114}: color_data = 12'h06b;
			{8'd86, 8'd115}: color_data = 12'h06b;
			{8'd86, 8'd116}: color_data = 12'h06b;
			{8'd86, 8'd117}: color_data = 12'h06b;
			{8'd86, 8'd118}: color_data = 12'h06b;
			{8'd86, 8'd119}: color_data = 12'h06b;
			{8'd86, 8'd120}: color_data = 12'h06b;
			{8'd86, 8'd121}: color_data = 12'h06b;
			{8'd86, 8'd122}: color_data = 12'h06b;
			{8'd86, 8'd123}: color_data = 12'h245;
			{8'd86, 8'd124}: color_data = 12'h432;
			{8'd86, 8'd125}: color_data = 12'h000;
			{8'd86, 8'd141}: color_data = 12'h000;
			{8'd86, 8'd142}: color_data = 12'h000;
			{8'd86, 8'd143}: color_data = 12'h210;
			{8'd86, 8'd144}: color_data = 12'h311;
			{8'd86, 8'd145}: color_data = 12'h210;
			{8'd86, 8'd146}: color_data = 12'h542;
			{8'd86, 8'd147}: color_data = 12'h964;
			{8'd86, 8'd148}: color_data = 12'h753;
			{8'd86, 8'd149}: color_data = 12'h000;
			{8'd87, 8'd7}: color_data = 12'hfc5;
			{8'd87, 8'd8}: color_data = 12'hfc3;
			{8'd87, 8'd9}: color_data = 12'hea0;
			{8'd87, 8'd10}: color_data = 12'hda0;
			{8'd87, 8'd11}: color_data = 12'hda0;
			{8'd87, 8'd12}: color_data = 12'heb3;
			{8'd87, 8'd13}: color_data = 12'hfc6;
			{8'd87, 8'd14}: color_data = 12'hfb3;
			{8'd87, 8'd15}: color_data = 12'hea0;
			{8'd87, 8'd16}: color_data = 12'hd90;
			{8'd87, 8'd17}: color_data = 12'heb2;
			{8'd87, 8'd18}: color_data = 12'hfc5;
			{8'd87, 8'd19}: color_data = 12'hd90;
			{8'd87, 8'd20}: color_data = 12'hd90;
			{8'd87, 8'd21}: color_data = 12'hd90;
			{8'd87, 8'd22}: color_data = 12'hea1;
			{8'd87, 8'd23}: color_data = 12'hfc5;
			{8'd87, 8'd24}: color_data = 12'hfc5;
			{8'd87, 8'd38}: color_data = 12'h000;
			{8'd87, 8'd39}: color_data = 12'h500;
			{8'd87, 8'd40}: color_data = 12'hd12;
			{8'd87, 8'd41}: color_data = 12'hf12;
			{8'd87, 8'd42}: color_data = 12'he12;
			{8'd87, 8'd43}: color_data = 12'he12;
			{8'd87, 8'd44}: color_data = 12'he12;
			{8'd87, 8'd45}: color_data = 12'he12;
			{8'd87, 8'd46}: color_data = 12'he12;
			{8'd87, 8'd47}: color_data = 12'he12;
			{8'd87, 8'd48}: color_data = 12'he12;
			{8'd87, 8'd49}: color_data = 12'he12;
			{8'd87, 8'd50}: color_data = 12'he12;
			{8'd87, 8'd51}: color_data = 12'he12;
			{8'd87, 8'd52}: color_data = 12'he12;
			{8'd87, 8'd53}: color_data = 12'he12;
			{8'd87, 8'd54}: color_data = 12'he12;
			{8'd87, 8'd55}: color_data = 12'he12;
			{8'd87, 8'd56}: color_data = 12'he12;
			{8'd87, 8'd57}: color_data = 12'he12;
			{8'd87, 8'd58}: color_data = 12'he12;
			{8'd87, 8'd59}: color_data = 12'hf12;
			{8'd87, 8'd60}: color_data = 12'hd12;
			{8'd87, 8'd61}: color_data = 12'h621;
			{8'd87, 8'd62}: color_data = 12'h843;
			{8'd87, 8'd63}: color_data = 12'h842;
			{8'd87, 8'd64}: color_data = 12'h842;
			{8'd87, 8'd65}: color_data = 12'h842;
			{8'd87, 8'd66}: color_data = 12'h843;
			{8'd87, 8'd67}: color_data = 12'h732;
			{8'd87, 8'd68}: color_data = 12'h976;
			{8'd87, 8'd69}: color_data = 12'hdb9;
			{8'd87, 8'd70}: color_data = 12'h986;
			{8'd87, 8'd71}: color_data = 12'heba;
			{8'd87, 8'd72}: color_data = 12'hfdb;
			{8'd87, 8'd73}: color_data = 12'hfda;
			{8'd87, 8'd74}: color_data = 12'hfda;
			{8'd87, 8'd75}: color_data = 12'hfda;
			{8'd87, 8'd76}: color_data = 12'hfdb;
			{8'd87, 8'd77}: color_data = 12'heca;
			{8'd87, 8'd78}: color_data = 12'h432;
			{8'd87, 8'd79}: color_data = 12'h976;
			{8'd87, 8'd80}: color_data = 12'h987;
			{8'd87, 8'd81}: color_data = 12'h059;
			{8'd87, 8'd82}: color_data = 12'h06b;
			{8'd87, 8'd83}: color_data = 12'h047;
			{8'd87, 8'd84}: color_data = 12'h612;
			{8'd87, 8'd85}: color_data = 12'hd11;
			{8'd87, 8'd86}: color_data = 12'hf12;
			{8'd87, 8'd87}: color_data = 12'hf12;
			{8'd87, 8'd88}: color_data = 12'he12;
			{8'd87, 8'd89}: color_data = 12'he12;
			{8'd87, 8'd90}: color_data = 12'he12;
			{8'd87, 8'd91}: color_data = 12'hf12;
			{8'd87, 8'd92}: color_data = 12'h912;
			{8'd87, 8'd93}: color_data = 12'h05a;
			{8'd87, 8'd94}: color_data = 12'h06b;
			{8'd87, 8'd95}: color_data = 12'h06b;
			{8'd87, 8'd96}: color_data = 12'h06b;
			{8'd87, 8'd97}: color_data = 12'h06b;
			{8'd87, 8'd98}: color_data = 12'h06b;
			{8'd87, 8'd99}: color_data = 12'h06b;
			{8'd87, 8'd100}: color_data = 12'h06b;
			{8'd87, 8'd101}: color_data = 12'h06b;
			{8'd87, 8'd102}: color_data = 12'h06b;
			{8'd87, 8'd103}: color_data = 12'h06b;
			{8'd87, 8'd104}: color_data = 12'h06b;
			{8'd87, 8'd105}: color_data = 12'h06b;
			{8'd87, 8'd106}: color_data = 12'h06b;
			{8'd87, 8'd107}: color_data = 12'h06b;
			{8'd87, 8'd108}: color_data = 12'h06b;
			{8'd87, 8'd109}: color_data = 12'h06b;
			{8'd87, 8'd110}: color_data = 12'h06b;
			{8'd87, 8'd111}: color_data = 12'h06b;
			{8'd87, 8'd112}: color_data = 12'h06b;
			{8'd87, 8'd113}: color_data = 12'h06b;
			{8'd87, 8'd114}: color_data = 12'h06b;
			{8'd87, 8'd115}: color_data = 12'h06b;
			{8'd87, 8'd116}: color_data = 12'h06b;
			{8'd87, 8'd117}: color_data = 12'h06b;
			{8'd87, 8'd118}: color_data = 12'h06b;
			{8'd87, 8'd119}: color_data = 12'h06b;
			{8'd87, 8'd120}: color_data = 12'h06b;
			{8'd87, 8'd121}: color_data = 12'h06b;
			{8'd87, 8'd122}: color_data = 12'h06b;
			{8'd87, 8'd123}: color_data = 12'h257;
			{8'd87, 8'd124}: color_data = 12'ha76;
			{8'd87, 8'd125}: color_data = 12'h322;
			{8'd87, 8'd140}: color_data = 12'h000;
			{8'd87, 8'd141}: color_data = 12'h311;
			{8'd87, 8'd142}: color_data = 12'h632;
			{8'd87, 8'd143}: color_data = 12'h842;
			{8'd87, 8'd144}: color_data = 12'h843;
			{8'd87, 8'd145}: color_data = 12'h842;
			{8'd87, 8'd146}: color_data = 12'h742;
			{8'd87, 8'd147}: color_data = 12'h753;
			{8'd87, 8'd148}: color_data = 12'hd95;
			{8'd87, 8'd149}: color_data = 12'hb84;
			{8'd87, 8'd150}: color_data = 12'h321;
			{8'd88, 8'd7}: color_data = 12'hfc4;
			{8'd88, 8'd8}: color_data = 12'hfd5;
			{8'd88, 8'd9}: color_data = 12'hfc5;
			{8'd88, 8'd10}: color_data = 12'hfc5;
			{8'd88, 8'd11}: color_data = 12'hfc5;
			{8'd88, 8'd12}: color_data = 12'hfc6;
			{8'd88, 8'd13}: color_data = 12'hfc5;
			{8'd88, 8'd14}: color_data = 12'hfc5;
			{8'd88, 8'd15}: color_data = 12'hfc5;
			{8'd88, 8'd16}: color_data = 12'hfc4;
			{8'd88, 8'd17}: color_data = 12'hfc6;
			{8'd88, 8'd18}: color_data = 12'hfc4;
			{8'd88, 8'd19}: color_data = 12'hd90;
			{8'd88, 8'd20}: color_data = 12'hd90;
			{8'd88, 8'd21}: color_data = 12'hd90;
			{8'd88, 8'd22}: color_data = 12'heb3;
			{8'd88, 8'd23}: color_data = 12'hfc5;
			{8'd88, 8'd24}: color_data = 12'hfc5;
			{8'd88, 8'd37}: color_data = 12'h000;
			{8'd88, 8'd38}: color_data = 12'h701;
			{8'd88, 8'd39}: color_data = 12'he12;
			{8'd88, 8'd40}: color_data = 12'hf12;
			{8'd88, 8'd41}: color_data = 12'he12;
			{8'd88, 8'd42}: color_data = 12'he12;
			{8'd88, 8'd43}: color_data = 12'he12;
			{8'd88, 8'd44}: color_data = 12'he12;
			{8'd88, 8'd45}: color_data = 12'he12;
			{8'd88, 8'd46}: color_data = 12'he12;
			{8'd88, 8'd47}: color_data = 12'he12;
			{8'd88, 8'd48}: color_data = 12'he12;
			{8'd88, 8'd49}: color_data = 12'he12;
			{8'd88, 8'd50}: color_data = 12'he12;
			{8'd88, 8'd51}: color_data = 12'he12;
			{8'd88, 8'd52}: color_data = 12'he12;
			{8'd88, 8'd53}: color_data = 12'he12;
			{8'd88, 8'd54}: color_data = 12'he12;
			{8'd88, 8'd55}: color_data = 12'he12;
			{8'd88, 8'd56}: color_data = 12'he12;
			{8'd88, 8'd57}: color_data = 12'he12;
			{8'd88, 8'd58}: color_data = 12'he12;
			{8'd88, 8'd59}: color_data = 12'he12;
			{8'd88, 8'd60}: color_data = 12'h711;
			{8'd88, 8'd61}: color_data = 12'h842;
			{8'd88, 8'd62}: color_data = 12'h842;
			{8'd88, 8'd63}: color_data = 12'h842;
			{8'd88, 8'd64}: color_data = 12'h842;
			{8'd88, 8'd65}: color_data = 12'h842;
			{8'd88, 8'd66}: color_data = 12'h842;
			{8'd88, 8'd67}: color_data = 12'h842;
			{8'd88, 8'd68}: color_data = 12'h632;
			{8'd88, 8'd69}: color_data = 12'hb97;
			{8'd88, 8'd70}: color_data = 12'heba;
			{8'd88, 8'd71}: color_data = 12'ha87;
			{8'd88, 8'd72}: color_data = 12'hda9;
			{8'd88, 8'd73}: color_data = 12'hfdb;
			{8'd88, 8'd74}: color_data = 12'hfda;
			{8'd88, 8'd75}: color_data = 12'hfda;
			{8'd88, 8'd76}: color_data = 12'hfdb;
			{8'd88, 8'd77}: color_data = 12'hb98;
			{8'd88, 8'd78}: color_data = 12'h865;
			{8'd88, 8'd79}: color_data = 12'hfdb;
			{8'd88, 8'd80}: color_data = 12'hfda;
			{8'd88, 8'd81}: color_data = 12'h456;
			{8'd88, 8'd82}: color_data = 12'h423;
			{8'd88, 8'd83}: color_data = 12'hc11;
			{8'd88, 8'd84}: color_data = 12'hf12;
			{8'd88, 8'd85}: color_data = 12'hf12;
			{8'd88, 8'd86}: color_data = 12'he12;
			{8'd88, 8'd87}: color_data = 12'he12;
			{8'd88, 8'd88}: color_data = 12'he12;
			{8'd88, 8'd89}: color_data = 12'he12;
			{8'd88, 8'd90}: color_data = 12'he12;
			{8'd88, 8'd91}: color_data = 12'hf12;
			{8'd88, 8'd92}: color_data = 12'ha12;
			{8'd88, 8'd93}: color_data = 12'h059;
			{8'd88, 8'd94}: color_data = 12'h06b;
			{8'd88, 8'd95}: color_data = 12'h06b;
			{8'd88, 8'd96}: color_data = 12'h06b;
			{8'd88, 8'd97}: color_data = 12'h06b;
			{8'd88, 8'd98}: color_data = 12'h06b;
			{8'd88, 8'd99}: color_data = 12'h06b;
			{8'd88, 8'd100}: color_data = 12'h06b;
			{8'd88, 8'd101}: color_data = 12'h06b;
			{8'd88, 8'd102}: color_data = 12'h06b;
			{8'd88, 8'd103}: color_data = 12'h06b;
			{8'd88, 8'd104}: color_data = 12'h06b;
			{8'd88, 8'd105}: color_data = 12'h06b;
			{8'd88, 8'd106}: color_data = 12'h06b;
			{8'd88, 8'd107}: color_data = 12'h06b;
			{8'd88, 8'd108}: color_data = 12'h06b;
			{8'd88, 8'd109}: color_data = 12'h06b;
			{8'd88, 8'd110}: color_data = 12'h06b;
			{8'd88, 8'd111}: color_data = 12'h06b;
			{8'd88, 8'd112}: color_data = 12'h06b;
			{8'd88, 8'd113}: color_data = 12'h06b;
			{8'd88, 8'd114}: color_data = 12'h06b;
			{8'd88, 8'd115}: color_data = 12'h06b;
			{8'd88, 8'd116}: color_data = 12'h06b;
			{8'd88, 8'd117}: color_data = 12'h06b;
			{8'd88, 8'd118}: color_data = 12'h06b;
			{8'd88, 8'd119}: color_data = 12'h06b;
			{8'd88, 8'd120}: color_data = 12'h06b;
			{8'd88, 8'd121}: color_data = 12'h06b;
			{8'd88, 8'd122}: color_data = 12'h06b;
			{8'd88, 8'd123}: color_data = 12'h047;
			{8'd88, 8'd124}: color_data = 12'hb86;
			{8'd88, 8'd125}: color_data = 12'h965;
			{8'd88, 8'd126}: color_data = 12'h000;
			{8'd88, 8'd139}: color_data = 12'h000;
			{8'd88, 8'd140}: color_data = 12'h421;
			{8'd88, 8'd141}: color_data = 12'h842;
			{8'd88, 8'd142}: color_data = 12'h843;
			{8'd88, 8'd143}: color_data = 12'h842;
			{8'd88, 8'd144}: color_data = 12'h842;
			{8'd88, 8'd145}: color_data = 12'h842;
			{8'd88, 8'd146}: color_data = 12'h843;
			{8'd88, 8'd147}: color_data = 12'h842;
			{8'd88, 8'd148}: color_data = 12'h632;
			{8'd88, 8'd149}: color_data = 12'hc95;
			{8'd88, 8'd150}: color_data = 12'hd95;
			{8'd88, 8'd151}: color_data = 12'h321;
			{8'd89, 8'd7}: color_data = 12'hfc5;
			{8'd89, 8'd8}: color_data = 12'hfc5;
			{8'd89, 8'd9}: color_data = 12'hfc5;
			{8'd89, 8'd10}: color_data = 12'hfc5;
			{8'd89, 8'd11}: color_data = 12'hfc5;
			{8'd89, 8'd12}: color_data = 12'hfc5;
			{8'd89, 8'd13}: color_data = 12'hfc6;
			{8'd89, 8'd14}: color_data = 12'hfc5;
			{8'd89, 8'd15}: color_data = 12'hfc5;
			{8'd89, 8'd16}: color_data = 12'hfc5;
			{8'd89, 8'd17}: color_data = 12'hfc5;
			{8'd89, 8'd18}: color_data = 12'hfc4;
			{8'd89, 8'd19}: color_data = 12'hd90;
			{8'd89, 8'd20}: color_data = 12'hd90;
			{8'd89, 8'd21}: color_data = 12'hd90;
			{8'd89, 8'd22}: color_data = 12'hfb3;
			{8'd89, 8'd23}: color_data = 12'hfc5;
			{8'd89, 8'd24}: color_data = 12'hfc5;
			{8'd89, 8'd36}: color_data = 12'h000;
			{8'd89, 8'd37}: color_data = 12'h701;
			{8'd89, 8'd38}: color_data = 12'hf12;
			{8'd89, 8'd39}: color_data = 12'hf12;
			{8'd89, 8'd40}: color_data = 12'he12;
			{8'd89, 8'd41}: color_data = 12'he12;
			{8'd89, 8'd42}: color_data = 12'he12;
			{8'd89, 8'd43}: color_data = 12'he12;
			{8'd89, 8'd44}: color_data = 12'he12;
			{8'd89, 8'd45}: color_data = 12'he12;
			{8'd89, 8'd46}: color_data = 12'he12;
			{8'd89, 8'd47}: color_data = 12'he12;
			{8'd89, 8'd48}: color_data = 12'he12;
			{8'd89, 8'd49}: color_data = 12'he12;
			{8'd89, 8'd50}: color_data = 12'he12;
			{8'd89, 8'd51}: color_data = 12'he12;
			{8'd89, 8'd52}: color_data = 12'he12;
			{8'd89, 8'd53}: color_data = 12'he12;
			{8'd89, 8'd54}: color_data = 12'he12;
			{8'd89, 8'd55}: color_data = 12'he12;
			{8'd89, 8'd56}: color_data = 12'he12;
			{8'd89, 8'd57}: color_data = 12'he12;
			{8'd89, 8'd58}: color_data = 12'hf12;
			{8'd89, 8'd59}: color_data = 12'h911;
			{8'd89, 8'd60}: color_data = 12'h742;
			{8'd89, 8'd61}: color_data = 12'h842;
			{8'd89, 8'd62}: color_data = 12'h643;
			{8'd89, 8'd63}: color_data = 12'h865;
			{8'd89, 8'd64}: color_data = 12'h632;
			{8'd89, 8'd65}: color_data = 12'h842;
			{8'd89, 8'd66}: color_data = 12'h842;
			{8'd89, 8'd67}: color_data = 12'h842;
			{8'd89, 8'd68}: color_data = 12'h842;
			{8'd89, 8'd69}: color_data = 12'h532;
			{8'd89, 8'd70}: color_data = 12'h765;
			{8'd89, 8'd71}: color_data = 12'hca8;
			{8'd89, 8'd72}: color_data = 12'hfca;
			{8'd89, 8'd73}: color_data = 12'hfdb;
			{8'd89, 8'd74}: color_data = 12'hfda;
			{8'd89, 8'd75}: color_data = 12'hfda;
			{8'd89, 8'd76}: color_data = 12'hfdb;
			{8'd89, 8'd77}: color_data = 12'hdb9;
			{8'd89, 8'd78}: color_data = 12'hfca;
			{8'd89, 8'd79}: color_data = 12'hfdb;
			{8'd89, 8'd80}: color_data = 12'hfdb;
			{8'd89, 8'd81}: color_data = 12'hb97;
			{8'd89, 8'd82}: color_data = 12'hc11;
			{8'd89, 8'd83}: color_data = 12'hf12;
			{8'd89, 8'd84}: color_data = 12'he12;
			{8'd89, 8'd85}: color_data = 12'he12;
			{8'd89, 8'd86}: color_data = 12'he12;
			{8'd89, 8'd87}: color_data = 12'he12;
			{8'd89, 8'd88}: color_data = 12'he12;
			{8'd89, 8'd89}: color_data = 12'he12;
			{8'd89, 8'd90}: color_data = 12'he12;
			{8'd89, 8'd91}: color_data = 12'hf12;
			{8'd89, 8'd92}: color_data = 12'hb11;
			{8'd89, 8'd93}: color_data = 12'h048;
			{8'd89, 8'd94}: color_data = 12'h06b;
			{8'd89, 8'd95}: color_data = 12'h06b;
			{8'd89, 8'd96}: color_data = 12'h06b;
			{8'd89, 8'd97}: color_data = 12'h06b;
			{8'd89, 8'd98}: color_data = 12'h06b;
			{8'd89, 8'd99}: color_data = 12'h06b;
			{8'd89, 8'd100}: color_data = 12'h06b;
			{8'd89, 8'd101}: color_data = 12'h06b;
			{8'd89, 8'd102}: color_data = 12'h06b;
			{8'd89, 8'd103}: color_data = 12'h06b;
			{8'd89, 8'd104}: color_data = 12'h06b;
			{8'd89, 8'd105}: color_data = 12'h06b;
			{8'd89, 8'd106}: color_data = 12'h06b;
			{8'd89, 8'd107}: color_data = 12'h06b;
			{8'd89, 8'd108}: color_data = 12'h06b;
			{8'd89, 8'd109}: color_data = 12'h06b;
			{8'd89, 8'd110}: color_data = 12'h06b;
			{8'd89, 8'd111}: color_data = 12'h06b;
			{8'd89, 8'd112}: color_data = 12'h06b;
			{8'd89, 8'd113}: color_data = 12'h06b;
			{8'd89, 8'd114}: color_data = 12'h06b;
			{8'd89, 8'd115}: color_data = 12'h06b;
			{8'd89, 8'd116}: color_data = 12'h06b;
			{8'd89, 8'd117}: color_data = 12'h06b;
			{8'd89, 8'd118}: color_data = 12'h06b;
			{8'd89, 8'd119}: color_data = 12'h06b;
			{8'd89, 8'd120}: color_data = 12'h06b;
			{8'd89, 8'd121}: color_data = 12'h06b;
			{8'd89, 8'd122}: color_data = 12'h06b;
			{8'd89, 8'd123}: color_data = 12'h058;
			{8'd89, 8'd124}: color_data = 12'h976;
			{8'd89, 8'd125}: color_data = 12'hc97;
			{8'd89, 8'd126}: color_data = 12'h432;
			{8'd89, 8'd139}: color_data = 12'h100;
			{8'd89, 8'd140}: color_data = 12'h742;
			{8'd89, 8'd141}: color_data = 12'h843;
			{8'd89, 8'd142}: color_data = 12'h842;
			{8'd89, 8'd143}: color_data = 12'h842;
			{8'd89, 8'd144}: color_data = 12'h842;
			{8'd89, 8'd145}: color_data = 12'h842;
			{8'd89, 8'd146}: color_data = 12'h842;
			{8'd89, 8'd147}: color_data = 12'h842;
			{8'd89, 8'd148}: color_data = 12'h842;
			{8'd89, 8'd149}: color_data = 12'h632;
			{8'd89, 8'd150}: color_data = 12'hd95;
			{8'd89, 8'd151}: color_data = 12'hc85;
			{8'd89, 8'd152}: color_data = 12'h110;
			{8'd90, 8'd8}: color_data = 12'hcc3;
			{8'd90, 8'd9}: color_data = 12'hec4;
			{8'd90, 8'd10}: color_data = 12'hec5;
			{8'd90, 8'd11}: color_data = 12'hec5;
			{8'd90, 8'd12}: color_data = 12'hfb5;
			{8'd90, 8'd14}: color_data = 12'hff0;
			{8'd90, 8'd15}: color_data = 12'hfd6;
			{8'd90, 8'd16}: color_data = 12'hfc5;
			{8'd90, 8'd17}: color_data = 12'hfc4;
			{8'd90, 8'd18}: color_data = 12'hfc5;
			{8'd90, 8'd19}: color_data = 12'hfc4;
			{8'd90, 8'd20}: color_data = 12'hea1;
			{8'd90, 8'd21}: color_data = 12'hd90;
			{8'd90, 8'd22}: color_data = 12'hfc4;
			{8'd90, 8'd23}: color_data = 12'hfc5;
			{8'd90, 8'd24}: color_data = 12'hfc5;
			{8'd90, 8'd35}: color_data = 12'h000;
			{8'd90, 8'd36}: color_data = 12'h701;
			{8'd90, 8'd37}: color_data = 12'hf12;
			{8'd90, 8'd38}: color_data = 12'hf12;
			{8'd90, 8'd39}: color_data = 12'he12;
			{8'd90, 8'd40}: color_data = 12'he12;
			{8'd90, 8'd41}: color_data = 12'he12;
			{8'd90, 8'd42}: color_data = 12'he12;
			{8'd90, 8'd43}: color_data = 12'he12;
			{8'd90, 8'd44}: color_data = 12'he12;
			{8'd90, 8'd45}: color_data = 12'he12;
			{8'd90, 8'd46}: color_data = 12'he12;
			{8'd90, 8'd47}: color_data = 12'he12;
			{8'd90, 8'd48}: color_data = 12'he12;
			{8'd90, 8'd49}: color_data = 12'he12;
			{8'd90, 8'd50}: color_data = 12'he12;
			{8'd90, 8'd51}: color_data = 12'he12;
			{8'd90, 8'd52}: color_data = 12'he12;
			{8'd90, 8'd53}: color_data = 12'he12;
			{8'd90, 8'd54}: color_data = 12'he12;
			{8'd90, 8'd55}: color_data = 12'he12;
			{8'd90, 8'd56}: color_data = 12'he12;
			{8'd90, 8'd57}: color_data = 12'hf12;
			{8'd90, 8'd58}: color_data = 12'hb11;
			{8'd90, 8'd59}: color_data = 12'h632;
			{8'd90, 8'd60}: color_data = 12'h842;
			{8'd90, 8'd61}: color_data = 12'h643;
			{8'd90, 8'd62}: color_data = 12'hdb9;
			{8'd90, 8'd63}: color_data = 12'hfdb;
			{8'd90, 8'd64}: color_data = 12'h875;
			{8'd90, 8'd65}: color_data = 12'h742;
			{8'd90, 8'd66}: color_data = 12'h843;
			{8'd90, 8'd67}: color_data = 12'h842;
			{8'd90, 8'd68}: color_data = 12'h842;
			{8'd90, 8'd69}: color_data = 12'h842;
			{8'd90, 8'd70}: color_data = 12'h643;
			{8'd90, 8'd71}: color_data = 12'hca8;
			{8'd90, 8'd72}: color_data = 12'heca;
			{8'd90, 8'd73}: color_data = 12'hfdb;
			{8'd90, 8'd74}: color_data = 12'hfda;
			{8'd90, 8'd75}: color_data = 12'hfda;
			{8'd90, 8'd76}: color_data = 12'hfda;
			{8'd90, 8'd77}: color_data = 12'hfdb;
			{8'd90, 8'd78}: color_data = 12'hfdb;
			{8'd90, 8'd79}: color_data = 12'hfda;
			{8'd90, 8'd80}: color_data = 12'hfdb;
			{8'd90, 8'd81}: color_data = 12'heca;
			{8'd90, 8'd82}: color_data = 12'h922;
			{8'd90, 8'd83}: color_data = 12'hf12;
			{8'd90, 8'd84}: color_data = 12'he12;
			{8'd90, 8'd85}: color_data = 12'he12;
			{8'd90, 8'd86}: color_data = 12'he12;
			{8'd90, 8'd87}: color_data = 12'he12;
			{8'd90, 8'd88}: color_data = 12'he12;
			{8'd90, 8'd89}: color_data = 12'he12;
			{8'd90, 8'd90}: color_data = 12'he12;
			{8'd90, 8'd91}: color_data = 12'hf12;
			{8'd90, 8'd92}: color_data = 12'hd11;
			{8'd90, 8'd93}: color_data = 12'h047;
			{8'd90, 8'd94}: color_data = 12'h06b;
			{8'd90, 8'd95}: color_data = 12'h06b;
			{8'd90, 8'd96}: color_data = 12'h06b;
			{8'd90, 8'd97}: color_data = 12'h06b;
			{8'd90, 8'd98}: color_data = 12'h06b;
			{8'd90, 8'd99}: color_data = 12'h06b;
			{8'd90, 8'd100}: color_data = 12'h06b;
			{8'd90, 8'd101}: color_data = 12'h06b;
			{8'd90, 8'd102}: color_data = 12'h06b;
			{8'd90, 8'd103}: color_data = 12'h06b;
			{8'd90, 8'd104}: color_data = 12'h06b;
			{8'd90, 8'd105}: color_data = 12'h06b;
			{8'd90, 8'd106}: color_data = 12'h06b;
			{8'd90, 8'd107}: color_data = 12'h06b;
			{8'd90, 8'd108}: color_data = 12'h06b;
			{8'd90, 8'd109}: color_data = 12'h06b;
			{8'd90, 8'd110}: color_data = 12'h06b;
			{8'd90, 8'd111}: color_data = 12'h06b;
			{8'd90, 8'd112}: color_data = 12'h06b;
			{8'd90, 8'd113}: color_data = 12'h06b;
			{8'd90, 8'd114}: color_data = 12'h06b;
			{8'd90, 8'd115}: color_data = 12'h06b;
			{8'd90, 8'd116}: color_data = 12'h06b;
			{8'd90, 8'd117}: color_data = 12'h06b;
			{8'd90, 8'd118}: color_data = 12'h06b;
			{8'd90, 8'd119}: color_data = 12'h06b;
			{8'd90, 8'd120}: color_data = 12'h06b;
			{8'd90, 8'd121}: color_data = 12'h06b;
			{8'd90, 8'd122}: color_data = 12'h06b;
			{8'd90, 8'd123}: color_data = 12'h059;
			{8'd90, 8'd124}: color_data = 12'h865;
			{8'd90, 8'd125}: color_data = 12'hda8;
			{8'd90, 8'd126}: color_data = 12'h864;
			{8'd90, 8'd127}: color_data = 12'h000;
			{8'd90, 8'd139}: color_data = 12'h321;
			{8'd90, 8'd140}: color_data = 12'h953;
			{8'd90, 8'd141}: color_data = 12'h843;
			{8'd90, 8'd142}: color_data = 12'h842;
			{8'd90, 8'd143}: color_data = 12'h842;
			{8'd90, 8'd144}: color_data = 12'h842;
			{8'd90, 8'd145}: color_data = 12'h842;
			{8'd90, 8'd146}: color_data = 12'h842;
			{8'd90, 8'd147}: color_data = 12'h842;
			{8'd90, 8'd148}: color_data = 12'h842;
			{8'd90, 8'd149}: color_data = 12'h842;
			{8'd90, 8'd150}: color_data = 12'h632;
			{8'd90, 8'd151}: color_data = 12'hea6;
			{8'd90, 8'd152}: color_data = 12'h863;
			{8'd91, 8'd17}: color_data = 12'hfc4;
			{8'd91, 8'd18}: color_data = 12'hfc5;
			{8'd91, 8'd19}: color_data = 12'hfc5;
			{8'd91, 8'd20}: color_data = 12'hfc5;
			{8'd91, 8'd21}: color_data = 12'hfb3;
			{8'd91, 8'd22}: color_data = 12'hfc5;
			{8'd91, 8'd23}: color_data = 12'hfc5;
			{8'd91, 8'd24}: color_data = 12'hfc6;
			{8'd91, 8'd34}: color_data = 12'h000;
			{8'd91, 8'd35}: color_data = 12'h701;
			{8'd91, 8'd36}: color_data = 12'hf12;
			{8'd91, 8'd37}: color_data = 12'hf12;
			{8'd91, 8'd38}: color_data = 12'he12;
			{8'd91, 8'd39}: color_data = 12'he12;
			{8'd91, 8'd40}: color_data = 12'he12;
			{8'd91, 8'd41}: color_data = 12'he12;
			{8'd91, 8'd42}: color_data = 12'he12;
			{8'd91, 8'd43}: color_data = 12'he12;
			{8'd91, 8'd44}: color_data = 12'he12;
			{8'd91, 8'd45}: color_data = 12'he12;
			{8'd91, 8'd46}: color_data = 12'he12;
			{8'd91, 8'd47}: color_data = 12'he12;
			{8'd91, 8'd48}: color_data = 12'he12;
			{8'd91, 8'd49}: color_data = 12'he12;
			{8'd91, 8'd50}: color_data = 12'he12;
			{8'd91, 8'd51}: color_data = 12'he12;
			{8'd91, 8'd52}: color_data = 12'he12;
			{8'd91, 8'd53}: color_data = 12'he12;
			{8'd91, 8'd54}: color_data = 12'he12;
			{8'd91, 8'd55}: color_data = 12'he12;
			{8'd91, 8'd56}: color_data = 12'hf12;
			{8'd91, 8'd57}: color_data = 12'hd12;
			{8'd91, 8'd58}: color_data = 12'h521;
			{8'd91, 8'd59}: color_data = 12'h732;
			{8'd91, 8'd60}: color_data = 12'h643;
			{8'd91, 8'd61}: color_data = 12'heb9;
			{8'd91, 8'd62}: color_data = 12'hfdb;
			{8'd91, 8'd63}: color_data = 12'hfdb;
			{8'd91, 8'd64}: color_data = 12'hdb9;
			{8'd91, 8'd65}: color_data = 12'h632;
			{8'd91, 8'd66}: color_data = 12'h842;
			{8'd91, 8'd67}: color_data = 12'h842;
			{8'd91, 8'd68}: color_data = 12'h842;
			{8'd91, 8'd69}: color_data = 12'h842;
			{8'd91, 8'd70}: color_data = 12'h643;
			{8'd91, 8'd71}: color_data = 12'heca;
			{8'd91, 8'd72}: color_data = 12'hfdb;
			{8'd91, 8'd73}: color_data = 12'hfda;
			{8'd91, 8'd74}: color_data = 12'hfda;
			{8'd91, 8'd75}: color_data = 12'hfda;
			{8'd91, 8'd76}: color_data = 12'hfda;
			{8'd91, 8'd77}: color_data = 12'hfda;
			{8'd91, 8'd78}: color_data = 12'hfda;
			{8'd91, 8'd79}: color_data = 12'hfda;
			{8'd91, 8'd80}: color_data = 12'hfda;
			{8'd91, 8'd81}: color_data = 12'hfdb;
			{8'd91, 8'd82}: color_data = 12'h944;
			{8'd91, 8'd83}: color_data = 12'he12;
			{8'd91, 8'd84}: color_data = 12'he12;
			{8'd91, 8'd85}: color_data = 12'he12;
			{8'd91, 8'd86}: color_data = 12'he12;
			{8'd91, 8'd87}: color_data = 12'he12;
			{8'd91, 8'd88}: color_data = 12'he12;
			{8'd91, 8'd89}: color_data = 12'he12;
			{8'd91, 8'd90}: color_data = 12'he12;
			{8'd91, 8'd91}: color_data = 12'he12;
			{8'd91, 8'd92}: color_data = 12'he11;
			{8'd91, 8'd93}: color_data = 12'h235;
			{8'd91, 8'd94}: color_data = 12'h06b;
			{8'd91, 8'd95}: color_data = 12'h06b;
			{8'd91, 8'd96}: color_data = 12'h06b;
			{8'd91, 8'd97}: color_data = 12'h06b;
			{8'd91, 8'd98}: color_data = 12'h06b;
			{8'd91, 8'd99}: color_data = 12'h06b;
			{8'd91, 8'd100}: color_data = 12'h06b;
			{8'd91, 8'd101}: color_data = 12'h06b;
			{8'd91, 8'd102}: color_data = 12'h06b;
			{8'd91, 8'd103}: color_data = 12'h06b;
			{8'd91, 8'd104}: color_data = 12'h06b;
			{8'd91, 8'd105}: color_data = 12'h06b;
			{8'd91, 8'd106}: color_data = 12'h06b;
			{8'd91, 8'd107}: color_data = 12'h06b;
			{8'd91, 8'd108}: color_data = 12'h06b;
			{8'd91, 8'd109}: color_data = 12'h06b;
			{8'd91, 8'd110}: color_data = 12'h06b;
			{8'd91, 8'd111}: color_data = 12'h06b;
			{8'd91, 8'd112}: color_data = 12'h06b;
			{8'd91, 8'd113}: color_data = 12'h06b;
			{8'd91, 8'd114}: color_data = 12'h06b;
			{8'd91, 8'd115}: color_data = 12'h06b;
			{8'd91, 8'd116}: color_data = 12'h06b;
			{8'd91, 8'd117}: color_data = 12'h06b;
			{8'd91, 8'd118}: color_data = 12'h06b;
			{8'd91, 8'd119}: color_data = 12'h06b;
			{8'd91, 8'd120}: color_data = 12'h06b;
			{8'd91, 8'd121}: color_data = 12'h06b;
			{8'd91, 8'd122}: color_data = 12'h06b;
			{8'd91, 8'd123}: color_data = 12'h05a;
			{8'd91, 8'd124}: color_data = 12'h655;
			{8'd91, 8'd125}: color_data = 12'hd97;
			{8'd91, 8'd126}: color_data = 12'ha86;
			{8'd91, 8'd127}: color_data = 12'h110;
			{8'd91, 8'd138}: color_data = 12'h000;
			{8'd91, 8'd139}: color_data = 12'h211;
			{8'd91, 8'd140}: color_data = 12'h632;
			{8'd91, 8'd141}: color_data = 12'h742;
			{8'd91, 8'd142}: color_data = 12'h842;
			{8'd91, 8'd143}: color_data = 12'h843;
			{8'd91, 8'd144}: color_data = 12'h842;
			{8'd91, 8'd145}: color_data = 12'h842;
			{8'd91, 8'd146}: color_data = 12'h842;
			{8'd91, 8'd147}: color_data = 12'h842;
			{8'd91, 8'd148}: color_data = 12'h842;
			{8'd91, 8'd149}: color_data = 12'h842;
			{8'd91, 8'd150}: color_data = 12'h842;
			{8'd91, 8'd151}: color_data = 12'h642;
			{8'd91, 8'd152}: color_data = 12'h642;
			{8'd91, 8'd153}: color_data = 12'h000;
			{8'd92, 8'd18}: color_data = 12'hfc4;
			{8'd92, 8'd19}: color_data = 12'hfc5;
			{8'd92, 8'd20}: color_data = 12'hfc5;
			{8'd92, 8'd21}: color_data = 12'hfc5;
			{8'd92, 8'd22}: color_data = 12'hfc4;
			{8'd92, 8'd23}: color_data = 12'hfc5;
			{8'd92, 8'd33}: color_data = 12'h000;
			{8'd92, 8'd34}: color_data = 12'h600;
			{8'd92, 8'd35}: color_data = 12'he12;
			{8'd92, 8'd36}: color_data = 12'hf12;
			{8'd92, 8'd37}: color_data = 12'he12;
			{8'd92, 8'd38}: color_data = 12'he12;
			{8'd92, 8'd39}: color_data = 12'he12;
			{8'd92, 8'd40}: color_data = 12'he12;
			{8'd92, 8'd41}: color_data = 12'he12;
			{8'd92, 8'd42}: color_data = 12'he12;
			{8'd92, 8'd43}: color_data = 12'he12;
			{8'd92, 8'd44}: color_data = 12'he12;
			{8'd92, 8'd45}: color_data = 12'he12;
			{8'd92, 8'd46}: color_data = 12'he12;
			{8'd92, 8'd47}: color_data = 12'he12;
			{8'd92, 8'd48}: color_data = 12'he12;
			{8'd92, 8'd49}: color_data = 12'he12;
			{8'd92, 8'd50}: color_data = 12'he12;
			{8'd92, 8'd51}: color_data = 12'he12;
			{8'd92, 8'd52}: color_data = 12'he12;
			{8'd92, 8'd53}: color_data = 12'he12;
			{8'd92, 8'd54}: color_data = 12'he12;
			{8'd92, 8'd55}: color_data = 12'he12;
			{8'd92, 8'd56}: color_data = 12'hf12;
			{8'd92, 8'd57}: color_data = 12'h801;
			{8'd92, 8'd58}: color_data = 12'h521;
			{8'd92, 8'd59}: color_data = 12'h976;
			{8'd92, 8'd60}: color_data = 12'hfca;
			{8'd92, 8'd61}: color_data = 12'hfdb;
			{8'd92, 8'd62}: color_data = 12'hfda;
			{8'd92, 8'd63}: color_data = 12'hfda;
			{8'd92, 8'd64}: color_data = 12'hfdb;
			{8'd92, 8'd65}: color_data = 12'h865;
			{8'd92, 8'd66}: color_data = 12'h742;
			{8'd92, 8'd67}: color_data = 12'h842;
			{8'd92, 8'd68}: color_data = 12'h842;
			{8'd92, 8'd69}: color_data = 12'h842;
			{8'd92, 8'd70}: color_data = 12'h643;
			{8'd92, 8'd71}: color_data = 12'hfca;
			{8'd92, 8'd72}: color_data = 12'hfdb;
			{8'd92, 8'd73}: color_data = 12'hfda;
			{8'd92, 8'd74}: color_data = 12'hfda;
			{8'd92, 8'd75}: color_data = 12'hfda;
			{8'd92, 8'd76}: color_data = 12'hfda;
			{8'd92, 8'd77}: color_data = 12'hfda;
			{8'd92, 8'd78}: color_data = 12'hfda;
			{8'd92, 8'd79}: color_data = 12'hfda;
			{8'd92, 8'd80}: color_data = 12'hfda;
			{8'd92, 8'd81}: color_data = 12'hfdb;
			{8'd92, 8'd82}: color_data = 12'ha65;
			{8'd92, 8'd83}: color_data = 12'he11;
			{8'd92, 8'd84}: color_data = 12'he12;
			{8'd92, 8'd85}: color_data = 12'he12;
			{8'd92, 8'd86}: color_data = 12'he12;
			{8'd92, 8'd87}: color_data = 12'he12;
			{8'd92, 8'd88}: color_data = 12'he12;
			{8'd92, 8'd89}: color_data = 12'he12;
			{8'd92, 8'd90}: color_data = 12'he12;
			{8'd92, 8'd91}: color_data = 12'he12;
			{8'd92, 8'd92}: color_data = 12'hf12;
			{8'd92, 8'd93}: color_data = 12'h623;
			{8'd92, 8'd94}: color_data = 12'h06b;
			{8'd92, 8'd95}: color_data = 12'h06b;
			{8'd92, 8'd96}: color_data = 12'h06b;
			{8'd92, 8'd97}: color_data = 12'h06b;
			{8'd92, 8'd98}: color_data = 12'h06b;
			{8'd92, 8'd99}: color_data = 12'h06b;
			{8'd92, 8'd100}: color_data = 12'h06b;
			{8'd92, 8'd101}: color_data = 12'h06b;
			{8'd92, 8'd102}: color_data = 12'h06b;
			{8'd92, 8'd103}: color_data = 12'h06b;
			{8'd92, 8'd104}: color_data = 12'h06b;
			{8'd92, 8'd105}: color_data = 12'h06b;
			{8'd92, 8'd106}: color_data = 12'h06b;
			{8'd92, 8'd107}: color_data = 12'h06b;
			{8'd92, 8'd108}: color_data = 12'h06b;
			{8'd92, 8'd109}: color_data = 12'h06b;
			{8'd92, 8'd110}: color_data = 12'h06b;
			{8'd92, 8'd111}: color_data = 12'h06b;
			{8'd92, 8'd112}: color_data = 12'h06b;
			{8'd92, 8'd113}: color_data = 12'h06b;
			{8'd92, 8'd114}: color_data = 12'h06b;
			{8'd92, 8'd115}: color_data = 12'h06b;
			{8'd92, 8'd116}: color_data = 12'h06b;
			{8'd92, 8'd117}: color_data = 12'h06b;
			{8'd92, 8'd118}: color_data = 12'h06b;
			{8'd92, 8'd119}: color_data = 12'h06b;
			{8'd92, 8'd120}: color_data = 12'h06b;
			{8'd92, 8'd121}: color_data = 12'h06b;
			{8'd92, 8'd122}: color_data = 12'h06b;
			{8'd92, 8'd123}: color_data = 12'h06b;
			{8'd92, 8'd124}: color_data = 12'h445;
			{8'd92, 8'd125}: color_data = 12'hd97;
			{8'd92, 8'd126}: color_data = 12'hc97;
			{8'd92, 8'd127}: color_data = 12'h432;
			{8'd92, 8'd137}: color_data = 12'h001;
			{8'd92, 8'd138}: color_data = 12'h035;
			{8'd92, 8'd139}: color_data = 12'h059;
			{8'd92, 8'd140}: color_data = 12'h059;
			{8'd92, 8'd141}: color_data = 12'h046;
			{8'd92, 8'd142}: color_data = 12'h433;
			{8'd92, 8'd143}: color_data = 12'h842;
			{8'd92, 8'd144}: color_data = 12'h843;
			{8'd92, 8'd145}: color_data = 12'h842;
			{8'd92, 8'd146}: color_data = 12'h842;
			{8'd92, 8'd147}: color_data = 12'h842;
			{8'd92, 8'd148}: color_data = 12'h842;
			{8'd92, 8'd149}: color_data = 12'h842;
			{8'd92, 8'd150}: color_data = 12'h843;
			{8'd92, 8'd151}: color_data = 12'h742;
			{8'd92, 8'd152}: color_data = 12'h753;
			{8'd92, 8'd153}: color_data = 12'h642;
			{8'd93, 8'd19}: color_data = 12'hff7;
			{8'd93, 8'd20}: color_data = 12'hfc5;
			{8'd93, 8'd21}: color_data = 12'hfc4;
			{8'd93, 8'd22}: color_data = 12'hfc4;
			{8'd93, 8'd23}: color_data = 12'hfd5;
			{8'd93, 8'd33}: color_data = 12'h400;
			{8'd93, 8'd34}: color_data = 12'hd12;
			{8'd93, 8'd35}: color_data = 12'hf12;
			{8'd93, 8'd36}: color_data = 12'he12;
			{8'd93, 8'd37}: color_data = 12'he12;
			{8'd93, 8'd38}: color_data = 12'he12;
			{8'd93, 8'd39}: color_data = 12'he12;
			{8'd93, 8'd40}: color_data = 12'he12;
			{8'd93, 8'd41}: color_data = 12'he12;
			{8'd93, 8'd42}: color_data = 12'he12;
			{8'd93, 8'd43}: color_data = 12'he12;
			{8'd93, 8'd44}: color_data = 12'he12;
			{8'd93, 8'd45}: color_data = 12'he12;
			{8'd93, 8'd46}: color_data = 12'he12;
			{8'd93, 8'd47}: color_data = 12'he12;
			{8'd93, 8'd48}: color_data = 12'he12;
			{8'd93, 8'd49}: color_data = 12'he12;
			{8'd93, 8'd50}: color_data = 12'he12;
			{8'd93, 8'd51}: color_data = 12'he12;
			{8'd93, 8'd52}: color_data = 12'he12;
			{8'd93, 8'd53}: color_data = 12'he12;
			{8'd93, 8'd54}: color_data = 12'he12;
			{8'd93, 8'd55}: color_data = 12'hf12;
			{8'd93, 8'd56}: color_data = 12'ha11;
			{8'd93, 8'd57}: color_data = 12'hb11;
			{8'd93, 8'd58}: color_data = 12'ha33;
			{8'd93, 8'd59}: color_data = 12'hfda;
			{8'd93, 8'd60}: color_data = 12'hfdb;
			{8'd93, 8'd61}: color_data = 12'hfda;
			{8'd93, 8'd62}: color_data = 12'hfda;
			{8'd93, 8'd63}: color_data = 12'hfda;
			{8'd93, 8'd64}: color_data = 12'hfdb;
			{8'd93, 8'd65}: color_data = 12'hca8;
			{8'd93, 8'd66}: color_data = 12'h632;
			{8'd93, 8'd67}: color_data = 12'h943;
			{8'd93, 8'd68}: color_data = 12'h632;
			{8'd93, 8'd69}: color_data = 12'h643;
			{8'd93, 8'd70}: color_data = 12'h976;
			{8'd93, 8'd71}: color_data = 12'hfdb;
			{8'd93, 8'd72}: color_data = 12'hfdb;
			{8'd93, 8'd73}: color_data = 12'hfda;
			{8'd93, 8'd74}: color_data = 12'hfda;
			{8'd93, 8'd75}: color_data = 12'hfda;
			{8'd93, 8'd76}: color_data = 12'hfda;
			{8'd93, 8'd77}: color_data = 12'hfda;
			{8'd93, 8'd78}: color_data = 12'hfda;
			{8'd93, 8'd79}: color_data = 12'hfda;
			{8'd93, 8'd80}: color_data = 12'hfda;
			{8'd93, 8'd81}: color_data = 12'hfdb;
			{8'd93, 8'd82}: color_data = 12'ha76;
			{8'd93, 8'd83}: color_data = 12'hd11;
			{8'd93, 8'd84}: color_data = 12'hf12;
			{8'd93, 8'd85}: color_data = 12'he12;
			{8'd93, 8'd86}: color_data = 12'he12;
			{8'd93, 8'd87}: color_data = 12'he12;
			{8'd93, 8'd88}: color_data = 12'hf12;
			{8'd93, 8'd89}: color_data = 12'hf12;
			{8'd93, 8'd90}: color_data = 12'hf12;
			{8'd93, 8'd91}: color_data = 12'hf12;
			{8'd93, 8'd92}: color_data = 12'hf11;
			{8'd93, 8'd93}: color_data = 12'h911;
			{8'd93, 8'd94}: color_data = 12'h048;
			{8'd93, 8'd95}: color_data = 12'h059;
			{8'd93, 8'd96}: color_data = 12'h058;
			{8'd93, 8'd97}: color_data = 12'h058;
			{8'd93, 8'd98}: color_data = 12'h059;
			{8'd93, 8'd99}: color_data = 12'h059;
			{8'd93, 8'd100}: color_data = 12'h06b;
			{8'd93, 8'd101}: color_data = 12'h06b;
			{8'd93, 8'd102}: color_data = 12'h06b;
			{8'd93, 8'd103}: color_data = 12'h06b;
			{8'd93, 8'd104}: color_data = 12'h06b;
			{8'd93, 8'd105}: color_data = 12'h06b;
			{8'd93, 8'd106}: color_data = 12'h06b;
			{8'd93, 8'd107}: color_data = 12'h06b;
			{8'd93, 8'd108}: color_data = 12'h06b;
			{8'd93, 8'd109}: color_data = 12'h06b;
			{8'd93, 8'd110}: color_data = 12'h06b;
			{8'd93, 8'd111}: color_data = 12'h06b;
			{8'd93, 8'd112}: color_data = 12'h06b;
			{8'd93, 8'd113}: color_data = 12'h06b;
			{8'd93, 8'd114}: color_data = 12'h06b;
			{8'd93, 8'd115}: color_data = 12'h06b;
			{8'd93, 8'd116}: color_data = 12'h06b;
			{8'd93, 8'd117}: color_data = 12'h06b;
			{8'd93, 8'd118}: color_data = 12'h06b;
			{8'd93, 8'd119}: color_data = 12'h06b;
			{8'd93, 8'd120}: color_data = 12'h06b;
			{8'd93, 8'd121}: color_data = 12'h06b;
			{8'd93, 8'd122}: color_data = 12'h06b;
			{8'd93, 8'd123}: color_data = 12'h06b;
			{8'd93, 8'd124}: color_data = 12'h059;
			{8'd93, 8'd125}: color_data = 12'h445;
			{8'd93, 8'd126}: color_data = 12'hb86;
			{8'd93, 8'd127}: color_data = 12'h754;
			{8'd93, 8'd136}: color_data = 12'h012;
			{8'd93, 8'd137}: color_data = 12'h048;
			{8'd93, 8'd138}: color_data = 12'h06b;
			{8'd93, 8'd139}: color_data = 12'h06b;
			{8'd93, 8'd140}: color_data = 12'h06b;
			{8'd93, 8'd141}: color_data = 12'h06b;
			{8'd93, 8'd142}: color_data = 12'h05a;
			{8'd93, 8'd143}: color_data = 12'h333;
			{8'd93, 8'd144}: color_data = 12'h842;
			{8'd93, 8'd145}: color_data = 12'h842;
			{8'd93, 8'd146}: color_data = 12'h842;
			{8'd93, 8'd147}: color_data = 12'h842;
			{8'd93, 8'd148}: color_data = 12'h842;
			{8'd93, 8'd149}: color_data = 12'h842;
			{8'd93, 8'd150}: color_data = 12'h842;
			{8'd93, 8'd151}: color_data = 12'h843;
			{8'd93, 8'd152}: color_data = 12'h632;
			{8'd93, 8'd153}: color_data = 12'h974;
			{8'd93, 8'd154}: color_data = 12'h431;
			{8'd94, 8'd21}: color_data = 12'hff0;
			{8'd94, 8'd32}: color_data = 12'h100;
			{8'd94, 8'd33}: color_data = 12'hb11;
			{8'd94, 8'd34}: color_data = 12'hf12;
			{8'd94, 8'd35}: color_data = 12'he12;
			{8'd94, 8'd36}: color_data = 12'he12;
			{8'd94, 8'd37}: color_data = 12'he12;
			{8'd94, 8'd38}: color_data = 12'he12;
			{8'd94, 8'd39}: color_data = 12'he12;
			{8'd94, 8'd40}: color_data = 12'he12;
			{8'd94, 8'd41}: color_data = 12'he12;
			{8'd94, 8'd42}: color_data = 12'he12;
			{8'd94, 8'd43}: color_data = 12'he12;
			{8'd94, 8'd44}: color_data = 12'he12;
			{8'd94, 8'd45}: color_data = 12'he12;
			{8'd94, 8'd46}: color_data = 12'he12;
			{8'd94, 8'd47}: color_data = 12'he12;
			{8'd94, 8'd48}: color_data = 12'he12;
			{8'd94, 8'd49}: color_data = 12'he12;
			{8'd94, 8'd50}: color_data = 12'he12;
			{8'd94, 8'd51}: color_data = 12'he12;
			{8'd94, 8'd52}: color_data = 12'he12;
			{8'd94, 8'd53}: color_data = 12'he12;
			{8'd94, 8'd54}: color_data = 12'hf12;
			{8'd94, 8'd55}: color_data = 12'hd12;
			{8'd94, 8'd56}: color_data = 12'h911;
			{8'd94, 8'd57}: color_data = 12'hf12;
			{8'd94, 8'd58}: color_data = 12'ha22;
			{8'd94, 8'd59}: color_data = 12'heca;
			{8'd94, 8'd60}: color_data = 12'hfdb;
			{8'd94, 8'd61}: color_data = 12'hfda;
			{8'd94, 8'd62}: color_data = 12'hfda;
			{8'd94, 8'd63}: color_data = 12'hfda;
			{8'd94, 8'd64}: color_data = 12'hfda;
			{8'd94, 8'd65}: color_data = 12'hfdb;
			{8'd94, 8'd66}: color_data = 12'h754;
			{8'd94, 8'd67}: color_data = 12'h732;
			{8'd94, 8'd68}: color_data = 12'h643;
			{8'd94, 8'd69}: color_data = 12'hb98;
			{8'd94, 8'd70}: color_data = 12'hb98;
			{8'd94, 8'd71}: color_data = 12'hca8;
			{8'd94, 8'd72}: color_data = 12'hfca;
			{8'd94, 8'd73}: color_data = 12'hfdb;
			{8'd94, 8'd74}: color_data = 12'hfda;
			{8'd94, 8'd75}: color_data = 12'hfda;
			{8'd94, 8'd76}: color_data = 12'hfda;
			{8'd94, 8'd77}: color_data = 12'hfda;
			{8'd94, 8'd78}: color_data = 12'hfda;
			{8'd94, 8'd79}: color_data = 12'hfda;
			{8'd94, 8'd80}: color_data = 12'hfda;
			{8'd94, 8'd81}: color_data = 12'hfdb;
			{8'd94, 8'd82}: color_data = 12'hb87;
			{8'd94, 8'd83}: color_data = 12'hc11;
			{8'd94, 8'd84}: color_data = 12'hf12;
			{8'd94, 8'd85}: color_data = 12'hf12;
			{8'd94, 8'd86}: color_data = 12'hf12;
			{8'd94, 8'd87}: color_data = 12'hf12;
			{8'd94, 8'd88}: color_data = 12'hd11;
			{8'd94, 8'd89}: color_data = 12'ha12;
			{8'd94, 8'd90}: color_data = 12'h713;
			{8'd94, 8'd91}: color_data = 12'h424;
			{8'd94, 8'd92}: color_data = 12'h235;
			{8'd94, 8'd93}: color_data = 12'h147;
			{8'd94, 8'd94}: color_data = 12'h048;
			{8'd94, 8'd95}: color_data = 12'h048;
			{8'd94, 8'd96}: color_data = 12'h048;
			{8'd94, 8'd97}: color_data = 12'h049;
			{8'd94, 8'd98}: color_data = 12'h058;
			{8'd94, 8'd99}: color_data = 12'h047;
			{8'd94, 8'd100}: color_data = 12'h036;
			{8'd94, 8'd101}: color_data = 12'h058;
			{8'd94, 8'd102}: color_data = 12'h06b;
			{8'd94, 8'd103}: color_data = 12'h06b;
			{8'd94, 8'd104}: color_data = 12'h06b;
			{8'd94, 8'd105}: color_data = 12'h06b;
			{8'd94, 8'd106}: color_data = 12'h06b;
			{8'd94, 8'd107}: color_data = 12'h06b;
			{8'd94, 8'd108}: color_data = 12'h06b;
			{8'd94, 8'd109}: color_data = 12'h06b;
			{8'd94, 8'd110}: color_data = 12'h06b;
			{8'd94, 8'd111}: color_data = 12'h06b;
			{8'd94, 8'd112}: color_data = 12'h06b;
			{8'd94, 8'd113}: color_data = 12'h06b;
			{8'd94, 8'd114}: color_data = 12'h06b;
			{8'd94, 8'd115}: color_data = 12'h06b;
			{8'd94, 8'd116}: color_data = 12'h06b;
			{8'd94, 8'd117}: color_data = 12'h06b;
			{8'd94, 8'd118}: color_data = 12'h06b;
			{8'd94, 8'd119}: color_data = 12'h06b;
			{8'd94, 8'd120}: color_data = 12'h06b;
			{8'd94, 8'd121}: color_data = 12'h06b;
			{8'd94, 8'd122}: color_data = 12'h06b;
			{8'd94, 8'd123}: color_data = 12'h06b;
			{8'd94, 8'd124}: color_data = 12'h06b;
			{8'd94, 8'd125}: color_data = 12'h05a;
			{8'd94, 8'd126}: color_data = 12'h147;
			{8'd94, 8'd127}: color_data = 12'h333;
			{8'd94, 8'd128}: color_data = 12'h000;
			{8'd94, 8'd135}: color_data = 12'h000;
			{8'd94, 8'd136}: color_data = 12'h048;
			{8'd94, 8'd137}: color_data = 12'h06b;
			{8'd94, 8'd138}: color_data = 12'h06b;
			{8'd94, 8'd139}: color_data = 12'h06b;
			{8'd94, 8'd140}: color_data = 12'h06b;
			{8'd94, 8'd141}: color_data = 12'h06b;
			{8'd94, 8'd142}: color_data = 12'h06b;
			{8'd94, 8'd143}: color_data = 12'h059;
			{8'd94, 8'd144}: color_data = 12'h432;
			{8'd94, 8'd145}: color_data = 12'h842;
			{8'd94, 8'd146}: color_data = 12'h842;
			{8'd94, 8'd147}: color_data = 12'h842;
			{8'd94, 8'd148}: color_data = 12'h842;
			{8'd94, 8'd149}: color_data = 12'h842;
			{8'd94, 8'd150}: color_data = 12'h842;
			{8'd94, 8'd151}: color_data = 12'h842;
			{8'd94, 8'd152}: color_data = 12'h842;
			{8'd94, 8'd153}: color_data = 12'h742;
			{8'd94, 8'd154}: color_data = 12'h974;
			{8'd94, 8'd155}: color_data = 12'h000;
			{8'd95, 8'd31}: color_data = 12'h000;
			{8'd95, 8'd32}: color_data = 12'h811;
			{8'd95, 8'd33}: color_data = 12'hf12;
			{8'd95, 8'd34}: color_data = 12'he12;
			{8'd95, 8'd35}: color_data = 12'he12;
			{8'd95, 8'd36}: color_data = 12'he12;
			{8'd95, 8'd37}: color_data = 12'he12;
			{8'd95, 8'd38}: color_data = 12'he12;
			{8'd95, 8'd39}: color_data = 12'he12;
			{8'd95, 8'd40}: color_data = 12'he12;
			{8'd95, 8'd41}: color_data = 12'he12;
			{8'd95, 8'd42}: color_data = 12'he12;
			{8'd95, 8'd43}: color_data = 12'he12;
			{8'd95, 8'd44}: color_data = 12'he12;
			{8'd95, 8'd45}: color_data = 12'he12;
			{8'd95, 8'd46}: color_data = 12'he12;
			{8'd95, 8'd47}: color_data = 12'he12;
			{8'd95, 8'd48}: color_data = 12'he12;
			{8'd95, 8'd49}: color_data = 12'hf12;
			{8'd95, 8'd50}: color_data = 12'hf12;
			{8'd95, 8'd51}: color_data = 12'hf12;
			{8'd95, 8'd52}: color_data = 12'hf12;
			{8'd95, 8'd53}: color_data = 12'he12;
			{8'd95, 8'd54}: color_data = 12'he12;
			{8'd95, 8'd55}: color_data = 12'h811;
			{8'd95, 8'd56}: color_data = 12'he12;
			{8'd95, 8'd57}: color_data = 12'hf12;
			{8'd95, 8'd58}: color_data = 12'h943;
			{8'd95, 8'd59}: color_data = 12'hfdb;
			{8'd95, 8'd60}: color_data = 12'hfdb;
			{8'd95, 8'd61}: color_data = 12'hfdb;
			{8'd95, 8'd62}: color_data = 12'hfda;
			{8'd95, 8'd63}: color_data = 12'hfda;
			{8'd95, 8'd64}: color_data = 12'hfda;
			{8'd95, 8'd65}: color_data = 12'hfdb;
			{8'd95, 8'd66}: color_data = 12'heba;
			{8'd95, 8'd67}: color_data = 12'h654;
			{8'd95, 8'd68}: color_data = 12'h765;
			{8'd95, 8'd69}: color_data = 12'hda9;
			{8'd95, 8'd70}: color_data = 12'hdb9;
			{8'd95, 8'd71}: color_data = 12'hca8;
			{8'd95, 8'd72}: color_data = 12'heba;
			{8'd95, 8'd73}: color_data = 12'hfdb;
			{8'd95, 8'd74}: color_data = 12'hfda;
			{8'd95, 8'd75}: color_data = 12'hfda;
			{8'd95, 8'd76}: color_data = 12'hfda;
			{8'd95, 8'd77}: color_data = 12'hfda;
			{8'd95, 8'd78}: color_data = 12'hfda;
			{8'd95, 8'd79}: color_data = 12'hfda;
			{8'd95, 8'd80}: color_data = 12'hfda;
			{8'd95, 8'd81}: color_data = 12'hfdb;
			{8'd95, 8'd82}: color_data = 12'hc98;
			{8'd95, 8'd83}: color_data = 12'hc11;
			{8'd95, 8'd84}: color_data = 12'hf11;
			{8'd95, 8'd85}: color_data = 12'hc11;
			{8'd95, 8'd86}: color_data = 12'ha11;
			{8'd95, 8'd87}: color_data = 12'h512;
			{8'd95, 8'd88}: color_data = 12'h124;
			{8'd95, 8'd89}: color_data = 12'h356;
			{8'd95, 8'd90}: color_data = 12'h257;
			{8'd95, 8'd91}: color_data = 12'h059;
			{8'd95, 8'd92}: color_data = 12'h06b;
			{8'd95, 8'd93}: color_data = 12'h05a;
			{8'd95, 8'd94}: color_data = 12'h156;
			{8'd95, 8'd95}: color_data = 12'h782;
			{8'd95, 8'd96}: color_data = 12'h891;
			{8'd95, 8'd97}: color_data = 12'h364;
			{8'd95, 8'd98}: color_data = 12'h059;
			{8'd95, 8'd99}: color_data = 12'h06b;
			{8'd95, 8'd100}: color_data = 12'h06b;
			{8'd95, 8'd101}: color_data = 12'h047;
			{8'd95, 8'd102}: color_data = 12'h048;
			{8'd95, 8'd103}: color_data = 12'h06b;
			{8'd95, 8'd104}: color_data = 12'h06b;
			{8'd95, 8'd105}: color_data = 12'h06b;
			{8'd95, 8'd106}: color_data = 12'h06b;
			{8'd95, 8'd107}: color_data = 12'h06b;
			{8'd95, 8'd108}: color_data = 12'h06b;
			{8'd95, 8'd109}: color_data = 12'h06b;
			{8'd95, 8'd110}: color_data = 12'h06b;
			{8'd95, 8'd111}: color_data = 12'h06b;
			{8'd95, 8'd112}: color_data = 12'h06b;
			{8'd95, 8'd113}: color_data = 12'h06b;
			{8'd95, 8'd114}: color_data = 12'h06b;
			{8'd95, 8'd115}: color_data = 12'h06b;
			{8'd95, 8'd116}: color_data = 12'h06b;
			{8'd95, 8'd117}: color_data = 12'h06b;
			{8'd95, 8'd118}: color_data = 12'h06b;
			{8'd95, 8'd119}: color_data = 12'h06b;
			{8'd95, 8'd120}: color_data = 12'h06b;
			{8'd95, 8'd121}: color_data = 12'h06b;
			{8'd95, 8'd122}: color_data = 12'h06b;
			{8'd95, 8'd123}: color_data = 12'h06b;
			{8'd95, 8'd124}: color_data = 12'h06b;
			{8'd95, 8'd125}: color_data = 12'h06b;
			{8'd95, 8'd126}: color_data = 12'h06b;
			{8'd95, 8'd127}: color_data = 12'h059;
			{8'd95, 8'd128}: color_data = 12'h025;
			{8'd95, 8'd129}: color_data = 12'h000;
			{8'd95, 8'd130}: color_data = 12'h000;
			{8'd95, 8'd132}: color_data = 12'h000;
			{8'd95, 8'd133}: color_data = 12'h013;
			{8'd95, 8'd134}: color_data = 12'h012;
			{8'd95, 8'd135}: color_data = 12'h013;
			{8'd95, 8'd136}: color_data = 12'h06b;
			{8'd95, 8'd137}: color_data = 12'h06b;
			{8'd95, 8'd138}: color_data = 12'h06b;
			{8'd95, 8'd139}: color_data = 12'h06b;
			{8'd95, 8'd140}: color_data = 12'h06b;
			{8'd95, 8'd141}: color_data = 12'h06b;
			{8'd95, 8'd142}: color_data = 12'h06b;
			{8'd95, 8'd143}: color_data = 12'h06b;
			{8'd95, 8'd144}: color_data = 12'h047;
			{8'd95, 8'd145}: color_data = 12'h732;
			{8'd95, 8'd146}: color_data = 12'h843;
			{8'd95, 8'd147}: color_data = 12'h842;
			{8'd95, 8'd148}: color_data = 12'h842;
			{8'd95, 8'd149}: color_data = 12'h842;
			{8'd95, 8'd150}: color_data = 12'h842;
			{8'd95, 8'd151}: color_data = 12'h842;
			{8'd95, 8'd152}: color_data = 12'h843;
			{8'd95, 8'd153}: color_data = 12'h732;
			{8'd95, 8'd154}: color_data = 12'ha74;
			{8'd95, 8'd155}: color_data = 12'h753;
			{8'd96, 8'd9}: color_data = 12'hfff;
			{8'd96, 8'd10}: color_data = 12'hfff;
			{8'd96, 8'd11}: color_data = 12'hfff;
			{8'd96, 8'd12}: color_data = 12'hfff;
			{8'd96, 8'd13}: color_data = 12'hfff;
			{8'd96, 8'd31}: color_data = 12'h400;
			{8'd96, 8'd32}: color_data = 12'he12;
			{8'd96, 8'd33}: color_data = 12'hf12;
			{8'd96, 8'd34}: color_data = 12'he12;
			{8'd96, 8'd35}: color_data = 12'he12;
			{8'd96, 8'd36}: color_data = 12'he12;
			{8'd96, 8'd37}: color_data = 12'he12;
			{8'd96, 8'd38}: color_data = 12'he12;
			{8'd96, 8'd39}: color_data = 12'he12;
			{8'd96, 8'd40}: color_data = 12'he12;
			{8'd96, 8'd41}: color_data = 12'he12;
			{8'd96, 8'd42}: color_data = 12'he12;
			{8'd96, 8'd43}: color_data = 12'he12;
			{8'd96, 8'd44}: color_data = 12'he12;
			{8'd96, 8'd45}: color_data = 12'he12;
			{8'd96, 8'd46}: color_data = 12'he12;
			{8'd96, 8'd47}: color_data = 12'hf12;
			{8'd96, 8'd48}: color_data = 12'he11;
			{8'd96, 8'd49}: color_data = 12'hc11;
			{8'd96, 8'd50}: color_data = 12'hb22;
			{8'd96, 8'd51}: color_data = 12'hb12;
			{8'd96, 8'd52}: color_data = 12'hc11;
			{8'd96, 8'd53}: color_data = 12'he11;
			{8'd96, 8'd54}: color_data = 12'ha11;
			{8'd96, 8'd55}: color_data = 12'hb11;
			{8'd96, 8'd56}: color_data = 12'hf12;
			{8'd96, 8'd57}: color_data = 12'hd11;
			{8'd96, 8'd58}: color_data = 12'ha76;
			{8'd96, 8'd59}: color_data = 12'hfdb;
			{8'd96, 8'd60}: color_data = 12'hfca;
			{8'd96, 8'd61}: color_data = 12'hfca;
			{8'd96, 8'd62}: color_data = 12'hfdb;
			{8'd96, 8'd63}: color_data = 12'hfdb;
			{8'd96, 8'd64}: color_data = 12'hfda;
			{8'd96, 8'd65}: color_data = 12'hfda;
			{8'd96, 8'd66}: color_data = 12'hfdb;
			{8'd96, 8'd67}: color_data = 12'ha87;
			{8'd96, 8'd68}: color_data = 12'heca;
			{8'd96, 8'd69}: color_data = 12'hfdb;
			{8'd96, 8'd70}: color_data = 12'hfdb;
			{8'd96, 8'd71}: color_data = 12'hfdb;
			{8'd96, 8'd72}: color_data = 12'hfdb;
			{8'd96, 8'd73}: color_data = 12'hfda;
			{8'd96, 8'd74}: color_data = 12'hfda;
			{8'd96, 8'd75}: color_data = 12'hfda;
			{8'd96, 8'd76}: color_data = 12'hfda;
			{8'd96, 8'd77}: color_data = 12'hfda;
			{8'd96, 8'd78}: color_data = 12'hfda;
			{8'd96, 8'd79}: color_data = 12'hfda;
			{8'd96, 8'd80}: color_data = 12'hfda;
			{8'd96, 8'd81}: color_data = 12'hfdb;
			{8'd96, 8'd82}: color_data = 12'hda8;
			{8'd96, 8'd83}: color_data = 12'h901;
			{8'd96, 8'd84}: color_data = 12'h944;
			{8'd96, 8'd85}: color_data = 12'hbbb;
			{8'd96, 8'd86}: color_data = 12'hcdd;
			{8'd96, 8'd87}: color_data = 12'h788;
			{8'd96, 8'd88}: color_data = 12'h9aa;
			{8'd96, 8'd89}: color_data = 12'hfff;
			{8'd96, 8'd90}: color_data = 12'hfff;
			{8'd96, 8'd91}: color_data = 12'h789;
			{8'd96, 8'd92}: color_data = 12'h357;
			{8'd96, 8'd93}: color_data = 12'h789;
			{8'd96, 8'd94}: color_data = 12'h874;
			{8'd96, 8'd95}: color_data = 12'hdd0;
			{8'd96, 8'd96}: color_data = 12'hfe0;
			{8'd96, 8'd97}: color_data = 12'hfe0;
			{8'd96, 8'd98}: color_data = 12'h990;
			{8'd96, 8'd99}: color_data = 12'h058;
			{8'd96, 8'd100}: color_data = 12'h06b;
			{8'd96, 8'd101}: color_data = 12'h06b;
			{8'd96, 8'd102}: color_data = 12'h036;
			{8'd96, 8'd103}: color_data = 12'h06a;
			{8'd96, 8'd104}: color_data = 12'h06b;
			{8'd96, 8'd105}: color_data = 12'h06b;
			{8'd96, 8'd106}: color_data = 12'h06b;
			{8'd96, 8'd107}: color_data = 12'h06b;
			{8'd96, 8'd108}: color_data = 12'h06b;
			{8'd96, 8'd109}: color_data = 12'h06b;
			{8'd96, 8'd110}: color_data = 12'h06b;
			{8'd96, 8'd111}: color_data = 12'h06b;
			{8'd96, 8'd112}: color_data = 12'h06b;
			{8'd96, 8'd113}: color_data = 12'h06b;
			{8'd96, 8'd114}: color_data = 12'h06b;
			{8'd96, 8'd115}: color_data = 12'h06b;
			{8'd96, 8'd116}: color_data = 12'h06b;
			{8'd96, 8'd117}: color_data = 12'h06b;
			{8'd96, 8'd118}: color_data = 12'h06b;
			{8'd96, 8'd119}: color_data = 12'h06b;
			{8'd96, 8'd120}: color_data = 12'h06b;
			{8'd96, 8'd121}: color_data = 12'h06b;
			{8'd96, 8'd122}: color_data = 12'h06b;
			{8'd96, 8'd123}: color_data = 12'h06b;
			{8'd96, 8'd124}: color_data = 12'h06b;
			{8'd96, 8'd125}: color_data = 12'h06b;
			{8'd96, 8'd126}: color_data = 12'h06b;
			{8'd96, 8'd127}: color_data = 12'h06b;
			{8'd96, 8'd128}: color_data = 12'h06b;
			{8'd96, 8'd129}: color_data = 12'h059;
			{8'd96, 8'd130}: color_data = 12'h036;
			{8'd96, 8'd131}: color_data = 12'h024;
			{8'd96, 8'd132}: color_data = 12'h013;
			{8'd96, 8'd133}: color_data = 12'h047;
			{8'd96, 8'd134}: color_data = 12'h05a;
			{8'd96, 8'd135}: color_data = 12'h048;
			{8'd96, 8'd136}: color_data = 12'h05a;
			{8'd96, 8'd137}: color_data = 12'h06b;
			{8'd96, 8'd138}: color_data = 12'h06b;
			{8'd96, 8'd139}: color_data = 12'h06b;
			{8'd96, 8'd140}: color_data = 12'h06b;
			{8'd96, 8'd141}: color_data = 12'h06b;
			{8'd96, 8'd142}: color_data = 12'h06b;
			{8'd96, 8'd143}: color_data = 12'h06b;
			{8'd96, 8'd144}: color_data = 12'h06b;
			{8'd96, 8'd145}: color_data = 12'h333;
			{8'd96, 8'd146}: color_data = 12'h842;
			{8'd96, 8'd147}: color_data = 12'h842;
			{8'd96, 8'd148}: color_data = 12'h842;
			{8'd96, 8'd149}: color_data = 12'h842;
			{8'd96, 8'd150}: color_data = 12'h842;
			{8'd96, 8'd151}: color_data = 12'h842;
			{8'd96, 8'd152}: color_data = 12'h842;
			{8'd96, 8'd153}: color_data = 12'h842;
			{8'd96, 8'd154}: color_data = 12'h642;
			{8'd96, 8'd155}: color_data = 12'hb84;
			{8'd96, 8'd156}: color_data = 12'h211;
			{8'd97, 8'd7}: color_data = 12'hfc5;
			{8'd97, 8'd8}: color_data = 12'hfc5;
			{8'd97, 8'd9}: color_data = 12'hfc5;
			{8'd97, 8'd10}: color_data = 12'hfc5;
			{8'd97, 8'd11}: color_data = 12'hfc5;
			{8'd97, 8'd12}: color_data = 12'hfc5;
			{8'd97, 8'd13}: color_data = 12'hfc5;
			{8'd97, 8'd14}: color_data = 12'hfc4;
			{8'd97, 8'd15}: color_data = 12'hfc5;
			{8'd97, 8'd16}: color_data = 12'hff0;
			{8'd97, 8'd30}: color_data = 12'h000;
			{8'd97, 8'd31}: color_data = 12'h911;
			{8'd97, 8'd32}: color_data = 12'hf12;
			{8'd97, 8'd33}: color_data = 12'he12;
			{8'd97, 8'd34}: color_data = 12'he12;
			{8'd97, 8'd35}: color_data = 12'he12;
			{8'd97, 8'd36}: color_data = 12'he12;
			{8'd97, 8'd37}: color_data = 12'he12;
			{8'd97, 8'd38}: color_data = 12'he12;
			{8'd97, 8'd39}: color_data = 12'he12;
			{8'd97, 8'd40}: color_data = 12'he12;
			{8'd97, 8'd41}: color_data = 12'he12;
			{8'd97, 8'd42}: color_data = 12'he12;
			{8'd97, 8'd43}: color_data = 12'he12;
			{8'd97, 8'd44}: color_data = 12'he12;
			{8'd97, 8'd45}: color_data = 12'he12;
			{8'd97, 8'd46}: color_data = 12'hf12;
			{8'd97, 8'd47}: color_data = 12'hd11;
			{8'd97, 8'd48}: color_data = 12'h945;
			{8'd97, 8'd49}: color_data = 12'hcbb;
			{8'd97, 8'd50}: color_data = 12'hdee;
			{8'd97, 8'd51}: color_data = 12'hddd;
			{8'd97, 8'd52}: color_data = 12'hbaa;
			{8'd97, 8'd53}: color_data = 12'h855;
			{8'd97, 8'd54}: color_data = 12'h901;
			{8'd97, 8'd55}: color_data = 12'hf12;
			{8'd97, 8'd56}: color_data = 12'hf12;
			{8'd97, 8'd57}: color_data = 12'ha11;
			{8'd97, 8'd58}: color_data = 12'h544;
			{8'd97, 8'd59}: color_data = 12'h432;
			{8'd97, 8'd60}: color_data = 12'h111;
			{8'd97, 8'd61}: color_data = 12'h221;
			{8'd97, 8'd62}: color_data = 12'h654;
			{8'd97, 8'd63}: color_data = 12'hca8;
			{8'd97, 8'd64}: color_data = 12'hfda;
			{8'd97, 8'd65}: color_data = 12'hfda;
			{8'd97, 8'd66}: color_data = 12'hfdb;
			{8'd97, 8'd67}: color_data = 12'hb98;
			{8'd97, 8'd68}: color_data = 12'hca8;
			{8'd97, 8'd69}: color_data = 12'hfdb;
			{8'd97, 8'd70}: color_data = 12'hdb9;
			{8'd97, 8'd71}: color_data = 12'ha86;
			{8'd97, 8'd72}: color_data = 12'hfca;
			{8'd97, 8'd73}: color_data = 12'hfdb;
			{8'd97, 8'd74}: color_data = 12'hfda;
			{8'd97, 8'd75}: color_data = 12'hfda;
			{8'd97, 8'd76}: color_data = 12'hfda;
			{8'd97, 8'd77}: color_data = 12'hfda;
			{8'd97, 8'd78}: color_data = 12'hfda;
			{8'd97, 8'd79}: color_data = 12'hfda;
			{8'd97, 8'd80}: color_data = 12'hfda;
			{8'd97, 8'd81}: color_data = 12'hfdb;
			{8'd97, 8'd82}: color_data = 12'hca8;
			{8'd97, 8'd83}: color_data = 12'h877;
			{8'd97, 8'd84}: color_data = 12'hfff;
			{8'd97, 8'd85}: color_data = 12'hfff;
			{8'd97, 8'd86}: color_data = 12'hfff;
			{8'd97, 8'd87}: color_data = 12'haaa;
			{8'd97, 8'd88}: color_data = 12'hfff;
			{8'd97, 8'd89}: color_data = 12'hfff;
			{8'd97, 8'd90}: color_data = 12'hfff;
			{8'd97, 8'd91}: color_data = 12'hfff;
			{8'd97, 8'd92}: color_data = 12'hfee;
			{8'd97, 8'd93}: color_data = 12'hfff;
			{8'd97, 8'd94}: color_data = 12'hfff;
			{8'd97, 8'd95}: color_data = 12'haa9;
			{8'd97, 8'd96}: color_data = 12'haa8;
			{8'd97, 8'd97}: color_data = 12'ha93;
			{8'd97, 8'd98}: color_data = 12'hba0;
			{8'd97, 8'd99}: color_data = 12'h058;
			{8'd97, 8'd100}: color_data = 12'h06b;
			{8'd97, 8'd101}: color_data = 12'h06b;
			{8'd97, 8'd102}: color_data = 12'h047;
			{8'd97, 8'd103}: color_data = 12'h05a;
			{8'd97, 8'd104}: color_data = 12'h06b;
			{8'd97, 8'd105}: color_data = 12'h06b;
			{8'd97, 8'd106}: color_data = 12'h06b;
			{8'd97, 8'd107}: color_data = 12'h06b;
			{8'd97, 8'd108}: color_data = 12'h06b;
			{8'd97, 8'd109}: color_data = 12'h06b;
			{8'd97, 8'd110}: color_data = 12'h06b;
			{8'd97, 8'd111}: color_data = 12'h06b;
			{8'd97, 8'd112}: color_data = 12'h06b;
			{8'd97, 8'd113}: color_data = 12'h06b;
			{8'd97, 8'd114}: color_data = 12'h06b;
			{8'd97, 8'd115}: color_data = 12'h06b;
			{8'd97, 8'd116}: color_data = 12'h06b;
			{8'd97, 8'd117}: color_data = 12'h06b;
			{8'd97, 8'd118}: color_data = 12'h06b;
			{8'd97, 8'd119}: color_data = 12'h06b;
			{8'd97, 8'd120}: color_data = 12'h06b;
			{8'd97, 8'd121}: color_data = 12'h06b;
			{8'd97, 8'd122}: color_data = 12'h06b;
			{8'd97, 8'd123}: color_data = 12'h06b;
			{8'd97, 8'd124}: color_data = 12'h06b;
			{8'd97, 8'd125}: color_data = 12'h06b;
			{8'd97, 8'd126}: color_data = 12'h06b;
			{8'd97, 8'd127}: color_data = 12'h06b;
			{8'd97, 8'd128}: color_data = 12'h06b;
			{8'd97, 8'd129}: color_data = 12'h06b;
			{8'd97, 8'd130}: color_data = 12'h06b;
			{8'd97, 8'd131}: color_data = 12'h06b;
			{8'd97, 8'd132}: color_data = 12'h05a;
			{8'd97, 8'd133}: color_data = 12'h059;
			{8'd97, 8'd134}: color_data = 12'h05a;
			{8'd97, 8'd135}: color_data = 12'h06b;
			{8'd97, 8'd136}: color_data = 12'h06b;
			{8'd97, 8'd137}: color_data = 12'h06b;
			{8'd97, 8'd138}: color_data = 12'h06b;
			{8'd97, 8'd139}: color_data = 12'h06b;
			{8'd97, 8'd140}: color_data = 12'h06b;
			{8'd97, 8'd141}: color_data = 12'h06b;
			{8'd97, 8'd142}: color_data = 12'h06b;
			{8'd97, 8'd143}: color_data = 12'h06b;
			{8'd97, 8'd144}: color_data = 12'h06b;
			{8'd97, 8'd145}: color_data = 12'h048;
			{8'd97, 8'd146}: color_data = 12'h732;
			{8'd97, 8'd147}: color_data = 12'h843;
			{8'd97, 8'd148}: color_data = 12'h842;
			{8'd97, 8'd149}: color_data = 12'h842;
			{8'd97, 8'd150}: color_data = 12'h842;
			{8'd97, 8'd151}: color_data = 12'h842;
			{8'd97, 8'd152}: color_data = 12'h842;
			{8'd97, 8'd153}: color_data = 12'h843;
			{8'd97, 8'd154}: color_data = 12'h742;
			{8'd97, 8'd155}: color_data = 12'h964;
			{8'd97, 8'd156}: color_data = 12'h863;
			{8'd97, 8'd157}: color_data = 12'h000;
			{8'd98, 8'd6}: color_data = 12'hfc5;
			{8'd98, 8'd7}: color_data = 12'hfc5;
			{8'd98, 8'd8}: color_data = 12'hfc5;
			{8'd98, 8'd9}: color_data = 12'hfc5;
			{8'd98, 8'd10}: color_data = 12'hfc5;
			{8'd98, 8'd11}: color_data = 12'hfc5;
			{8'd98, 8'd12}: color_data = 12'hfc5;
			{8'd98, 8'd13}: color_data = 12'hfc5;
			{8'd98, 8'd14}: color_data = 12'hfc5;
			{8'd98, 8'd15}: color_data = 12'hfc5;
			{8'd98, 8'd16}: color_data = 12'hfc5;
			{8'd98, 8'd17}: color_data = 12'hfc6;
			{8'd98, 8'd30}: color_data = 12'h000;
			{8'd98, 8'd31}: color_data = 12'h911;
			{8'd98, 8'd32}: color_data = 12'hf12;
			{8'd98, 8'd33}: color_data = 12'he12;
			{8'd98, 8'd34}: color_data = 12'he12;
			{8'd98, 8'd35}: color_data = 12'he12;
			{8'd98, 8'd36}: color_data = 12'he12;
			{8'd98, 8'd37}: color_data = 12'he12;
			{8'd98, 8'd38}: color_data = 12'he12;
			{8'd98, 8'd39}: color_data = 12'he12;
			{8'd98, 8'd40}: color_data = 12'he12;
			{8'd98, 8'd41}: color_data = 12'he12;
			{8'd98, 8'd42}: color_data = 12'he12;
			{8'd98, 8'd43}: color_data = 12'he12;
			{8'd98, 8'd44}: color_data = 12'he12;
			{8'd98, 8'd45}: color_data = 12'hf12;
			{8'd98, 8'd46}: color_data = 12'hd11;
			{8'd98, 8'd47}: color_data = 12'h966;
			{8'd98, 8'd48}: color_data = 12'hfff;
			{8'd98, 8'd49}: color_data = 12'hfff;
			{8'd98, 8'd50}: color_data = 12'hfff;
			{8'd98, 8'd51}: color_data = 12'hfff;
			{8'd98, 8'd52}: color_data = 12'hfff;
			{8'd98, 8'd53}: color_data = 12'h977;
			{8'd98, 8'd54}: color_data = 12'hd11;
			{8'd98, 8'd55}: color_data = 12'hf12;
			{8'd98, 8'd56}: color_data = 12'hf12;
			{8'd98, 8'd57}: color_data = 12'h400;
			{8'd98, 8'd58}: color_data = 12'h000;
			{8'd98, 8'd59}: color_data = 12'h433;
			{8'd98, 8'd60}: color_data = 12'h865;
			{8'd98, 8'd61}: color_data = 12'ha87;
			{8'd98, 8'd62}: color_data = 12'h986;
			{8'd98, 8'd63}: color_data = 12'ha87;
			{8'd98, 8'd64}: color_data = 12'hfca;
			{8'd98, 8'd65}: color_data = 12'hfdb;
			{8'd98, 8'd66}: color_data = 12'hfdb;
			{8'd98, 8'd67}: color_data = 12'hfca;
			{8'd98, 8'd68}: color_data = 12'heba;
			{8'd98, 8'd69}: color_data = 12'hfdb;
			{8'd98, 8'd70}: color_data = 12'hfdb;
			{8'd98, 8'd71}: color_data = 12'hdb9;
			{8'd98, 8'd72}: color_data = 12'h976;
			{8'd98, 8'd73}: color_data = 12'hfda;
			{8'd98, 8'd74}: color_data = 12'hfdb;
			{8'd98, 8'd75}: color_data = 12'hfda;
			{8'd98, 8'd76}: color_data = 12'hfda;
			{8'd98, 8'd77}: color_data = 12'hfda;
			{8'd98, 8'd78}: color_data = 12'hfda;
			{8'd98, 8'd79}: color_data = 12'hfda;
			{8'd98, 8'd80}: color_data = 12'hfdb;
			{8'd98, 8'd81}: color_data = 12'hfca;
			{8'd98, 8'd82}: color_data = 12'h988;
			{8'd98, 8'd83}: color_data = 12'hfff;
			{8'd98, 8'd84}: color_data = 12'hfff;
			{8'd98, 8'd85}: color_data = 12'hfff;
			{8'd98, 8'd86}: color_data = 12'hfff;
			{8'd98, 8'd87}: color_data = 12'hddd;
			{8'd98, 8'd88}: color_data = 12'hfff;
			{8'd98, 8'd89}: color_data = 12'hfff;
			{8'd98, 8'd90}: color_data = 12'hfff;
			{8'd98, 8'd91}: color_data = 12'hfff;
			{8'd98, 8'd92}: color_data = 12'hfff;
			{8'd98, 8'd93}: color_data = 12'hfff;
			{8'd98, 8'd94}: color_data = 12'hfff;
			{8'd98, 8'd95}: color_data = 12'hfff;
			{8'd98, 8'd96}: color_data = 12'hfff;
			{8'd98, 8'd97}: color_data = 12'hedd;
			{8'd98, 8'd98}: color_data = 12'h135;
			{8'd98, 8'd99}: color_data = 12'h049;
			{8'd98, 8'd100}: color_data = 12'h059;
			{8'd98, 8'd101}: color_data = 12'h048;
			{8'd98, 8'd102}: color_data = 12'h047;
			{8'd98, 8'd103}: color_data = 12'h06b;
			{8'd98, 8'd104}: color_data = 12'h06b;
			{8'd98, 8'd105}: color_data = 12'h06b;
			{8'd98, 8'd106}: color_data = 12'h06b;
			{8'd98, 8'd107}: color_data = 12'h06b;
			{8'd98, 8'd108}: color_data = 12'h06b;
			{8'd98, 8'd109}: color_data = 12'h06b;
			{8'd98, 8'd110}: color_data = 12'h06b;
			{8'd98, 8'd111}: color_data = 12'h06b;
			{8'd98, 8'd112}: color_data = 12'h06b;
			{8'd98, 8'd113}: color_data = 12'h06b;
			{8'd98, 8'd114}: color_data = 12'h06b;
			{8'd98, 8'd115}: color_data = 12'h06b;
			{8'd98, 8'd116}: color_data = 12'h06b;
			{8'd98, 8'd117}: color_data = 12'h06b;
			{8'd98, 8'd118}: color_data = 12'h06b;
			{8'd98, 8'd119}: color_data = 12'h06b;
			{8'd98, 8'd120}: color_data = 12'h06b;
			{8'd98, 8'd121}: color_data = 12'h06b;
			{8'd98, 8'd122}: color_data = 12'h06b;
			{8'd98, 8'd123}: color_data = 12'h06b;
			{8'd98, 8'd124}: color_data = 12'h06b;
			{8'd98, 8'd125}: color_data = 12'h06b;
			{8'd98, 8'd126}: color_data = 12'h06b;
			{8'd98, 8'd127}: color_data = 12'h06b;
			{8'd98, 8'd128}: color_data = 12'h06b;
			{8'd98, 8'd129}: color_data = 12'h06b;
			{8'd98, 8'd130}: color_data = 12'h06b;
			{8'd98, 8'd131}: color_data = 12'h06b;
			{8'd98, 8'd132}: color_data = 12'h06b;
			{8'd98, 8'd133}: color_data = 12'h06b;
			{8'd98, 8'd134}: color_data = 12'h06b;
			{8'd98, 8'd135}: color_data = 12'h06b;
			{8'd98, 8'd136}: color_data = 12'h06b;
			{8'd98, 8'd137}: color_data = 12'h06b;
			{8'd98, 8'd138}: color_data = 12'h06b;
			{8'd98, 8'd139}: color_data = 12'h06b;
			{8'd98, 8'd140}: color_data = 12'h06b;
			{8'd98, 8'd141}: color_data = 12'h06b;
			{8'd98, 8'd142}: color_data = 12'h06b;
			{8'd98, 8'd143}: color_data = 12'h06b;
			{8'd98, 8'd144}: color_data = 12'h06b;
			{8'd98, 8'd145}: color_data = 12'h06a;
			{8'd98, 8'd146}: color_data = 12'h333;
			{8'd98, 8'd147}: color_data = 12'h842;
			{8'd98, 8'd148}: color_data = 12'h843;
			{8'd98, 8'd149}: color_data = 12'h842;
			{8'd98, 8'd150}: color_data = 12'h842;
			{8'd98, 8'd151}: color_data = 12'h842;
			{8'd98, 8'd152}: color_data = 12'h842;
			{8'd98, 8'd153}: color_data = 12'h842;
			{8'd98, 8'd154}: color_data = 12'h842;
			{8'd98, 8'd155}: color_data = 12'h642;
			{8'd98, 8'd156}: color_data = 12'ha74;
			{8'd98, 8'd157}: color_data = 12'h110;
			{8'd99, 8'd5}: color_data = 12'hfc5;
			{8'd99, 8'd6}: color_data = 12'hfc5;
			{8'd99, 8'd7}: color_data = 12'hfc5;
			{8'd99, 8'd8}: color_data = 12'hfb3;
			{8'd99, 8'd9}: color_data = 12'hea1;
			{8'd99, 8'd10}: color_data = 12'hea1;
			{8'd99, 8'd11}: color_data = 12'hea1;
			{8'd99, 8'd12}: color_data = 12'hea1;
			{8'd99, 8'd13}: color_data = 12'hea1;
			{8'd99, 8'd14}: color_data = 12'heb3;
			{8'd99, 8'd15}: color_data = 12'hfc5;
			{8'd99, 8'd16}: color_data = 12'hfc5;
			{8'd99, 8'd17}: color_data = 12'hfc5;
			{8'd99, 8'd18}: color_data = 12'heb5;
			{8'd99, 8'd31}: color_data = 12'h601;
			{8'd99, 8'd32}: color_data = 12'hf12;
			{8'd99, 8'd33}: color_data = 12'he12;
			{8'd99, 8'd34}: color_data = 12'he12;
			{8'd99, 8'd35}: color_data = 12'he12;
			{8'd99, 8'd36}: color_data = 12'he12;
			{8'd99, 8'd37}: color_data = 12'he12;
			{8'd99, 8'd38}: color_data = 12'he12;
			{8'd99, 8'd39}: color_data = 12'he12;
			{8'd99, 8'd40}: color_data = 12'he12;
			{8'd99, 8'd41}: color_data = 12'he12;
			{8'd99, 8'd42}: color_data = 12'he12;
			{8'd99, 8'd43}: color_data = 12'he12;
			{8'd99, 8'd44}: color_data = 12'he12;
			{8'd99, 8'd45}: color_data = 12'he12;
			{8'd99, 8'd46}: color_data = 12'h933;
			{8'd99, 8'd47}: color_data = 12'heff;
			{8'd99, 8'd48}: color_data = 12'hfff;
			{8'd99, 8'd49}: color_data = 12'hfff;
			{8'd99, 8'd50}: color_data = 12'hfee;
			{8'd99, 8'd51}: color_data = 12'hfee;
			{8'd99, 8'd52}: color_data = 12'hcbb;
			{8'd99, 8'd53}: color_data = 12'ha12;
			{8'd99, 8'd54}: color_data = 12'hf12;
			{8'd99, 8'd55}: color_data = 12'hf12;
			{8'd99, 8'd56}: color_data = 12'hc11;
			{8'd99, 8'd57}: color_data = 12'h876;
			{8'd99, 8'd58}: color_data = 12'heca;
			{8'd99, 8'd59}: color_data = 12'hfdb;
			{8'd99, 8'd60}: color_data = 12'hfdb;
			{8'd99, 8'd61}: color_data = 12'hfdb;
			{8'd99, 8'd62}: color_data = 12'hfdb;
			{8'd99, 8'd63}: color_data = 12'hfdb;
			{8'd99, 8'd64}: color_data = 12'hfda;
			{8'd99, 8'd65}: color_data = 12'hfda;
			{8'd99, 8'd66}: color_data = 12'hfdb;
			{8'd99, 8'd67}: color_data = 12'hfca;
			{8'd99, 8'd68}: color_data = 12'h543;
			{8'd99, 8'd69}: color_data = 12'h322;
			{8'd99, 8'd70}: color_data = 12'ha87;
			{8'd99, 8'd71}: color_data = 12'hfdb;
			{8'd99, 8'd72}: color_data = 12'hb98;
			{8'd99, 8'd73}: color_data = 12'h332;
			{8'd99, 8'd74}: color_data = 12'hdb9;
			{8'd99, 8'd75}: color_data = 12'hfdb;
			{8'd99, 8'd76}: color_data = 12'hfda;
			{8'd99, 8'd77}: color_data = 12'hfda;
			{8'd99, 8'd78}: color_data = 12'hfda;
			{8'd99, 8'd79}: color_data = 12'hfda;
			{8'd99, 8'd80}: color_data = 12'hfdb;
			{8'd99, 8'd81}: color_data = 12'hdb9;
			{8'd99, 8'd82}: color_data = 12'hbba;
			{8'd99, 8'd83}: color_data = 12'hfff;
			{8'd99, 8'd84}: color_data = 12'hfff;
			{8'd99, 8'd85}: color_data = 12'hfff;
			{8'd99, 8'd86}: color_data = 12'hfff;
			{8'd99, 8'd87}: color_data = 12'hfff;
			{8'd99, 8'd88}: color_data = 12'hfff;
			{8'd99, 8'd89}: color_data = 12'hfff;
			{8'd99, 8'd90}: color_data = 12'hfff;
			{8'd99, 8'd91}: color_data = 12'hfff;
			{8'd99, 8'd92}: color_data = 12'hfff;
			{8'd99, 8'd93}: color_data = 12'hfff;
			{8'd99, 8'd94}: color_data = 12'hfff;
			{8'd99, 8'd95}: color_data = 12'hfff;
			{8'd99, 8'd96}: color_data = 12'hfff;
			{8'd99, 8'd97}: color_data = 12'hccc;
			{8'd99, 8'd98}: color_data = 12'h765;
			{8'd99, 8'd99}: color_data = 12'h654;
			{8'd99, 8'd100}: color_data = 12'h134;
			{8'd99, 8'd101}: color_data = 12'h048;
			{8'd99, 8'd102}: color_data = 12'h06b;
			{8'd99, 8'd103}: color_data = 12'h06b;
			{8'd99, 8'd104}: color_data = 12'h06b;
			{8'd99, 8'd105}: color_data = 12'h06b;
			{8'd99, 8'd106}: color_data = 12'h06b;
			{8'd99, 8'd107}: color_data = 12'h06b;
			{8'd99, 8'd108}: color_data = 12'h06b;
			{8'd99, 8'd109}: color_data = 12'h06b;
			{8'd99, 8'd110}: color_data = 12'h06b;
			{8'd99, 8'd111}: color_data = 12'h06b;
			{8'd99, 8'd112}: color_data = 12'h06b;
			{8'd99, 8'd113}: color_data = 12'h06b;
			{8'd99, 8'd114}: color_data = 12'h06b;
			{8'd99, 8'd115}: color_data = 12'h06b;
			{8'd99, 8'd116}: color_data = 12'h06b;
			{8'd99, 8'd117}: color_data = 12'h06b;
			{8'd99, 8'd118}: color_data = 12'h06b;
			{8'd99, 8'd119}: color_data = 12'h06b;
			{8'd99, 8'd120}: color_data = 12'h06b;
			{8'd99, 8'd121}: color_data = 12'h06b;
			{8'd99, 8'd122}: color_data = 12'h06b;
			{8'd99, 8'd123}: color_data = 12'h06b;
			{8'd99, 8'd124}: color_data = 12'h06b;
			{8'd99, 8'd125}: color_data = 12'h06b;
			{8'd99, 8'd126}: color_data = 12'h06b;
			{8'd99, 8'd127}: color_data = 12'h06b;
			{8'd99, 8'd128}: color_data = 12'h06b;
			{8'd99, 8'd129}: color_data = 12'h06b;
			{8'd99, 8'd130}: color_data = 12'h06b;
			{8'd99, 8'd131}: color_data = 12'h06b;
			{8'd99, 8'd132}: color_data = 12'h06b;
			{8'd99, 8'd133}: color_data = 12'h06b;
			{8'd99, 8'd134}: color_data = 12'h06b;
			{8'd99, 8'd135}: color_data = 12'h06b;
			{8'd99, 8'd136}: color_data = 12'h06b;
			{8'd99, 8'd137}: color_data = 12'h06b;
			{8'd99, 8'd138}: color_data = 12'h06b;
			{8'd99, 8'd139}: color_data = 12'h06b;
			{8'd99, 8'd140}: color_data = 12'h06b;
			{8'd99, 8'd141}: color_data = 12'h06b;
			{8'd99, 8'd142}: color_data = 12'h06b;
			{8'd99, 8'd143}: color_data = 12'h06b;
			{8'd99, 8'd144}: color_data = 12'h06b;
			{8'd99, 8'd145}: color_data = 12'h06b;
			{8'd99, 8'd146}: color_data = 12'h136;
			{8'd99, 8'd147}: color_data = 12'h842;
			{8'd99, 8'd148}: color_data = 12'h742;
			{8'd99, 8'd149}: color_data = 12'h842;
			{8'd99, 8'd150}: color_data = 12'h842;
			{8'd99, 8'd151}: color_data = 12'h842;
			{8'd99, 8'd152}: color_data = 12'h842;
			{8'd99, 8'd153}: color_data = 12'h842;
			{8'd99, 8'd154}: color_data = 12'h843;
			{8'd99, 8'd155}: color_data = 12'h742;
			{8'd99, 8'd156}: color_data = 12'h964;
			{8'd99, 8'd157}: color_data = 12'h642;
			{8'd100, 8'd4}: color_data = 12'hfc5;
			{8'd100, 8'd5}: color_data = 12'hfc5;
			{8'd100, 8'd6}: color_data = 12'hfc5;
			{8'd100, 8'd7}: color_data = 12'hfb3;
			{8'd100, 8'd8}: color_data = 12'hd90;
			{8'd100, 8'd9}: color_data = 12'hd90;
			{8'd100, 8'd10}: color_data = 12'hd90;
			{8'd100, 8'd11}: color_data = 12'hd90;
			{8'd100, 8'd12}: color_data = 12'hd90;
			{8'd100, 8'd13}: color_data = 12'hd90;
			{8'd100, 8'd14}: color_data = 12'hd90;
			{8'd100, 8'd15}: color_data = 12'hea1;
			{8'd100, 8'd16}: color_data = 12'hfc4;
			{8'd100, 8'd17}: color_data = 12'hfc5;
			{8'd100, 8'd18}: color_data = 12'hfc5;
			{8'd100, 8'd19}: color_data = 12'hfc6;
			{8'd100, 8'd31}: color_data = 12'h300;
			{8'd100, 8'd32}: color_data = 12'hd12;
			{8'd100, 8'd33}: color_data = 12'hf12;
			{8'd100, 8'd34}: color_data = 12'he12;
			{8'd100, 8'd35}: color_data = 12'he12;
			{8'd100, 8'd36}: color_data = 12'he12;
			{8'd100, 8'd37}: color_data = 12'he12;
			{8'd100, 8'd38}: color_data = 12'he12;
			{8'd100, 8'd39}: color_data = 12'he12;
			{8'd100, 8'd40}: color_data = 12'he12;
			{8'd100, 8'd41}: color_data = 12'he12;
			{8'd100, 8'd42}: color_data = 12'he12;
			{8'd100, 8'd43}: color_data = 12'he12;
			{8'd100, 8'd44}: color_data = 12'hf12;
			{8'd100, 8'd45}: color_data = 12'hc11;
			{8'd100, 8'd46}: color_data = 12'hbaa;
			{8'd100, 8'd47}: color_data = 12'hfff;
			{8'd100, 8'd48}: color_data = 12'hf99;
			{8'd100, 8'd49}: color_data = 12'hfab;
			{8'd100, 8'd50}: color_data = 12'hfbb;
			{8'd100, 8'd51}: color_data = 12'hfcc;
			{8'd100, 8'd52}: color_data = 12'h933;
			{8'd100, 8'd53}: color_data = 12'he11;
			{8'd100, 8'd54}: color_data = 12'he12;
			{8'd100, 8'd55}: color_data = 12'he12;
			{8'd100, 8'd56}: color_data = 12'h943;
			{8'd100, 8'd57}: color_data = 12'hdb9;
			{8'd100, 8'd58}: color_data = 12'hb97;
			{8'd100, 8'd59}: color_data = 12'ha87;
			{8'd100, 8'd60}: color_data = 12'ha87;
			{8'd100, 8'd61}: color_data = 12'ha87;
			{8'd100, 8'd62}: color_data = 12'hb98;
			{8'd100, 8'd63}: color_data = 12'heb9;
			{8'd100, 8'd64}: color_data = 12'hfdb;
			{8'd100, 8'd65}: color_data = 12'hfda;
			{8'd100, 8'd66}: color_data = 12'hfda;
			{8'd100, 8'd67}: color_data = 12'hfdb;
			{8'd100, 8'd68}: color_data = 12'h765;
			{8'd100, 8'd69}: color_data = 12'h000;
			{8'd100, 8'd70}: color_data = 12'h000;
			{8'd100, 8'd71}: color_data = 12'h976;
			{8'd100, 8'd72}: color_data = 12'hca8;
			{8'd100, 8'd73}: color_data = 12'h000;
			{8'd100, 8'd74}: color_data = 12'h765;
			{8'd100, 8'd75}: color_data = 12'hfdb;
			{8'd100, 8'd76}: color_data = 12'hfda;
			{8'd100, 8'd77}: color_data = 12'hfda;
			{8'd100, 8'd78}: color_data = 12'hfda;
			{8'd100, 8'd79}: color_data = 12'hfda;
			{8'd100, 8'd80}: color_data = 12'hfdb;
			{8'd100, 8'd81}: color_data = 12'hdb9;
			{8'd100, 8'd82}: color_data = 12'hbbb;
			{8'd100, 8'd83}: color_data = 12'hfff;
			{8'd100, 8'd84}: color_data = 12'hfff;
			{8'd100, 8'd85}: color_data = 12'hfff;
			{8'd100, 8'd86}: color_data = 12'hfff;
			{8'd100, 8'd87}: color_data = 12'hfff;
			{8'd100, 8'd88}: color_data = 12'hfff;
			{8'd100, 8'd89}: color_data = 12'hfff;
			{8'd100, 8'd90}: color_data = 12'hfff;
			{8'd100, 8'd91}: color_data = 12'hfff;
			{8'd100, 8'd92}: color_data = 12'hfff;
			{8'd100, 8'd93}: color_data = 12'hfff;
			{8'd100, 8'd94}: color_data = 12'hfff;
			{8'd100, 8'd95}: color_data = 12'hfff;
			{8'd100, 8'd96}: color_data = 12'hfff;
			{8'd100, 8'd97}: color_data = 12'hbbb;
			{8'd100, 8'd98}: color_data = 12'h975;
			{8'd100, 8'd99}: color_data = 12'hda7;
			{8'd100, 8'd100}: color_data = 12'hb86;
			{8'd100, 8'd101}: color_data = 12'h655;
			{8'd100, 8'd102}: color_data = 12'h047;
			{8'd100, 8'd103}: color_data = 12'h05a;
			{8'd100, 8'd104}: color_data = 12'h06b;
			{8'd100, 8'd105}: color_data = 12'h06b;
			{8'd100, 8'd106}: color_data = 12'h06b;
			{8'd100, 8'd107}: color_data = 12'h06b;
			{8'd100, 8'd108}: color_data = 12'h06b;
			{8'd100, 8'd109}: color_data = 12'h06b;
			{8'd100, 8'd110}: color_data = 12'h06b;
			{8'd100, 8'd111}: color_data = 12'h06b;
			{8'd100, 8'd112}: color_data = 12'h06b;
			{8'd100, 8'd113}: color_data = 12'h06b;
			{8'd100, 8'd114}: color_data = 12'h06b;
			{8'd100, 8'd115}: color_data = 12'h06b;
			{8'd100, 8'd116}: color_data = 12'h06b;
			{8'd100, 8'd117}: color_data = 12'h06b;
			{8'd100, 8'd118}: color_data = 12'h06b;
			{8'd100, 8'd119}: color_data = 12'h06b;
			{8'd100, 8'd120}: color_data = 12'h06b;
			{8'd100, 8'd121}: color_data = 12'h06b;
			{8'd100, 8'd122}: color_data = 12'h06b;
			{8'd100, 8'd123}: color_data = 12'h06b;
			{8'd100, 8'd124}: color_data = 12'h06b;
			{8'd100, 8'd125}: color_data = 12'h06b;
			{8'd100, 8'd126}: color_data = 12'h06b;
			{8'd100, 8'd127}: color_data = 12'h06b;
			{8'd100, 8'd128}: color_data = 12'h06b;
			{8'd100, 8'd129}: color_data = 12'h06b;
			{8'd100, 8'd130}: color_data = 12'h06b;
			{8'd100, 8'd131}: color_data = 12'h06b;
			{8'd100, 8'd132}: color_data = 12'h06b;
			{8'd100, 8'd133}: color_data = 12'h06b;
			{8'd100, 8'd134}: color_data = 12'h06b;
			{8'd100, 8'd135}: color_data = 12'h06b;
			{8'd100, 8'd136}: color_data = 12'h06b;
			{8'd100, 8'd137}: color_data = 12'h06b;
			{8'd100, 8'd138}: color_data = 12'h06b;
			{8'd100, 8'd139}: color_data = 12'h06b;
			{8'd100, 8'd140}: color_data = 12'h06b;
			{8'd100, 8'd141}: color_data = 12'h06b;
			{8'd100, 8'd142}: color_data = 12'h06b;
			{8'd100, 8'd143}: color_data = 12'h06b;
			{8'd100, 8'd144}: color_data = 12'h06b;
			{8'd100, 8'd145}: color_data = 12'h06b;
			{8'd100, 8'd146}: color_data = 12'h048;
			{8'd100, 8'd147}: color_data = 12'h632;
			{8'd100, 8'd148}: color_data = 12'h531;
			{8'd100, 8'd149}: color_data = 12'h843;
			{8'd100, 8'd150}: color_data = 12'h842;
			{8'd100, 8'd151}: color_data = 12'h842;
			{8'd100, 8'd152}: color_data = 12'h842;
			{8'd100, 8'd153}: color_data = 12'h842;
			{8'd100, 8'd154}: color_data = 12'h842;
			{8'd100, 8'd155}: color_data = 12'h842;
			{8'd100, 8'd156}: color_data = 12'h742;
			{8'd100, 8'd157}: color_data = 12'h863;
			{8'd100, 8'd158}: color_data = 12'h000;
			{8'd101, 8'd3}: color_data = 12'hfc6;
			{8'd101, 8'd4}: color_data = 12'hfc5;
			{8'd101, 8'd5}: color_data = 12'hfc5;
			{8'd101, 8'd6}: color_data = 12'heb3;
			{8'd101, 8'd7}: color_data = 12'hd90;
			{8'd101, 8'd8}: color_data = 12'hd90;
			{8'd101, 8'd9}: color_data = 12'hd90;
			{8'd101, 8'd10}: color_data = 12'hd90;
			{8'd101, 8'd11}: color_data = 12'hd90;
			{8'd101, 8'd12}: color_data = 12'hd90;
			{8'd101, 8'd13}: color_data = 12'hd90;
			{8'd101, 8'd14}: color_data = 12'hd90;
			{8'd101, 8'd15}: color_data = 12'hd90;
			{8'd101, 8'd16}: color_data = 12'hda0;
			{8'd101, 8'd17}: color_data = 12'hfb3;
			{8'd101, 8'd18}: color_data = 12'hfc5;
			{8'd101, 8'd19}: color_data = 12'hfc5;
			{8'd101, 8'd20}: color_data = 12'hfc5;
			{8'd101, 8'd31}: color_data = 12'h000;
			{8'd101, 8'd32}: color_data = 12'h811;
			{8'd101, 8'd33}: color_data = 12'hf12;
			{8'd101, 8'd34}: color_data = 12'he12;
			{8'd101, 8'd35}: color_data = 12'he12;
			{8'd101, 8'd36}: color_data = 12'he12;
			{8'd101, 8'd37}: color_data = 12'he12;
			{8'd101, 8'd38}: color_data = 12'he12;
			{8'd101, 8'd39}: color_data = 12'he12;
			{8'd101, 8'd40}: color_data = 12'he12;
			{8'd101, 8'd41}: color_data = 12'he12;
			{8'd101, 8'd42}: color_data = 12'he12;
			{8'd101, 8'd43}: color_data = 12'he12;
			{8'd101, 8'd44}: color_data = 12'hf12;
			{8'd101, 8'd45}: color_data = 12'ha33;
			{8'd101, 8'd46}: color_data = 12'heff;
			{8'd101, 8'd47}: color_data = 12'hfff;
			{8'd101, 8'd48}: color_data = 12'hfcc;
			{8'd101, 8'd49}: color_data = 12'hfbb;
			{8'd101, 8'd50}: color_data = 12'hfff;
			{8'd101, 8'd51}: color_data = 12'hbbb;
			{8'd101, 8'd52}: color_data = 12'hc11;
			{8'd101, 8'd53}: color_data = 12'hf12;
			{8'd101, 8'd54}: color_data = 12'hf12;
			{8'd101, 8'd55}: color_data = 12'hb11;
			{8'd101, 8'd56}: color_data = 12'h654;
			{8'd101, 8'd57}: color_data = 12'hb97;
			{8'd101, 8'd58}: color_data = 12'heb9;
			{8'd101, 8'd59}: color_data = 12'hfca;
			{8'd101, 8'd60}: color_data = 12'hfca;
			{8'd101, 8'd61}: color_data = 12'heca;
			{8'd101, 8'd62}: color_data = 12'hca8;
			{8'd101, 8'd63}: color_data = 12'ha87;
			{8'd101, 8'd64}: color_data = 12'hca8;
			{8'd101, 8'd65}: color_data = 12'hfdb;
			{8'd101, 8'd66}: color_data = 12'hfdb;
			{8'd101, 8'd67}: color_data = 12'hfdb;
			{8'd101, 8'd68}: color_data = 12'heba;
			{8'd101, 8'd69}: color_data = 12'h111;
			{8'd101, 8'd70}: color_data = 12'h000;
			{8'd101, 8'd71}: color_data = 12'h000;
			{8'd101, 8'd72}: color_data = 12'h221;
			{8'd101, 8'd73}: color_data = 12'h000;
			{8'd101, 8'd74}: color_data = 12'h543;
			{8'd101, 8'd75}: color_data = 12'hfdb;
			{8'd101, 8'd76}: color_data = 12'hfda;
			{8'd101, 8'd77}: color_data = 12'hfda;
			{8'd101, 8'd78}: color_data = 12'hfda;
			{8'd101, 8'd79}: color_data = 12'hfda;
			{8'd101, 8'd80}: color_data = 12'hfdb;
			{8'd101, 8'd81}: color_data = 12'hdb9;
			{8'd101, 8'd82}: color_data = 12'h999;
			{8'd101, 8'd83}: color_data = 12'hfff;
			{8'd101, 8'd84}: color_data = 12'hfff;
			{8'd101, 8'd85}: color_data = 12'hfff;
			{8'd101, 8'd86}: color_data = 12'hfff;
			{8'd101, 8'd87}: color_data = 12'hfff;
			{8'd101, 8'd88}: color_data = 12'hfff;
			{8'd101, 8'd89}: color_data = 12'hfff;
			{8'd101, 8'd90}: color_data = 12'hfff;
			{8'd101, 8'd91}: color_data = 12'hfff;
			{8'd101, 8'd92}: color_data = 12'hfff;
			{8'd101, 8'd93}: color_data = 12'hfff;
			{8'd101, 8'd94}: color_data = 12'hfff;
			{8'd101, 8'd95}: color_data = 12'hfff;
			{8'd101, 8'd96}: color_data = 12'hfff;
			{8'd101, 8'd97}: color_data = 12'hfff;
			{8'd101, 8'd98}: color_data = 12'h876;
			{8'd101, 8'd99}: color_data = 12'hc97;
			{8'd101, 8'd100}: color_data = 12'hc97;
			{8'd101, 8'd101}: color_data = 12'hd97;
			{8'd101, 8'd102}: color_data = 12'ha86;
			{8'd101, 8'd103}: color_data = 12'h445;
			{8'd101, 8'd104}: color_data = 12'h059;
			{8'd101, 8'd105}: color_data = 12'h06b;
			{8'd101, 8'd106}: color_data = 12'h06b;
			{8'd101, 8'd107}: color_data = 12'h06b;
			{8'd101, 8'd108}: color_data = 12'h06b;
			{8'd101, 8'd109}: color_data = 12'h06b;
			{8'd101, 8'd110}: color_data = 12'h06b;
			{8'd101, 8'd111}: color_data = 12'h06b;
			{8'd101, 8'd112}: color_data = 12'h06b;
			{8'd101, 8'd113}: color_data = 12'h06b;
			{8'd101, 8'd114}: color_data = 12'h06b;
			{8'd101, 8'd115}: color_data = 12'h06b;
			{8'd101, 8'd116}: color_data = 12'h06b;
			{8'd101, 8'd117}: color_data = 12'h06b;
			{8'd101, 8'd118}: color_data = 12'h06b;
			{8'd101, 8'd119}: color_data = 12'h06b;
			{8'd101, 8'd120}: color_data = 12'h06b;
			{8'd101, 8'd121}: color_data = 12'h06b;
			{8'd101, 8'd122}: color_data = 12'h06b;
			{8'd101, 8'd123}: color_data = 12'h06b;
			{8'd101, 8'd124}: color_data = 12'h06b;
			{8'd101, 8'd125}: color_data = 12'h06b;
			{8'd101, 8'd126}: color_data = 12'h06b;
			{8'd101, 8'd127}: color_data = 12'h06b;
			{8'd101, 8'd128}: color_data = 12'h06b;
			{8'd101, 8'd129}: color_data = 12'h06b;
			{8'd101, 8'd130}: color_data = 12'h06b;
			{8'd101, 8'd131}: color_data = 12'h06b;
			{8'd101, 8'd132}: color_data = 12'h06b;
			{8'd101, 8'd133}: color_data = 12'h06b;
			{8'd101, 8'd134}: color_data = 12'h06b;
			{8'd101, 8'd135}: color_data = 12'h06b;
			{8'd101, 8'd136}: color_data = 12'h06b;
			{8'd101, 8'd137}: color_data = 12'h06b;
			{8'd101, 8'd138}: color_data = 12'h06b;
			{8'd101, 8'd139}: color_data = 12'h06b;
			{8'd101, 8'd140}: color_data = 12'h06b;
			{8'd101, 8'd141}: color_data = 12'h06b;
			{8'd101, 8'd142}: color_data = 12'h06b;
			{8'd101, 8'd143}: color_data = 12'h06b;
			{8'd101, 8'd144}: color_data = 12'h06b;
			{8'd101, 8'd145}: color_data = 12'h06b;
			{8'd101, 8'd146}: color_data = 12'h059;
			{8'd101, 8'd147}: color_data = 12'h321;
			{8'd101, 8'd148}: color_data = 12'h742;
			{8'd101, 8'd149}: color_data = 12'h843;
			{8'd101, 8'd150}: color_data = 12'h842;
			{8'd101, 8'd151}: color_data = 12'h842;
			{8'd101, 8'd152}: color_data = 12'h842;
			{8'd101, 8'd153}: color_data = 12'h842;
			{8'd101, 8'd154}: color_data = 12'h842;
			{8'd101, 8'd155}: color_data = 12'h843;
			{8'd101, 8'd156}: color_data = 12'h742;
			{8'd101, 8'd157}: color_data = 12'h863;
			{8'd101, 8'd158}: color_data = 12'h211;
			{8'd102, 8'd3}: color_data = 12'hfc5;
			{8'd102, 8'd4}: color_data = 12'hfc5;
			{8'd102, 8'd5}: color_data = 12'heb2;
			{8'd102, 8'd6}: color_data = 12'hd90;
			{8'd102, 8'd7}: color_data = 12'hd90;
			{8'd102, 8'd8}: color_data = 12'hd90;
			{8'd102, 8'd9}: color_data = 12'hd90;
			{8'd102, 8'd10}: color_data = 12'hd90;
			{8'd102, 8'd11}: color_data = 12'hd90;
			{8'd102, 8'd12}: color_data = 12'hd90;
			{8'd102, 8'd13}: color_data = 12'hd90;
			{8'd102, 8'd14}: color_data = 12'hd90;
			{8'd102, 8'd15}: color_data = 12'hd90;
			{8'd102, 8'd16}: color_data = 12'hd90;
			{8'd102, 8'd17}: color_data = 12'hd90;
			{8'd102, 8'd18}: color_data = 12'heb2;
			{8'd102, 8'd19}: color_data = 12'hfc5;
			{8'd102, 8'd20}: color_data = 12'hfc5;
			{8'd102, 8'd21}: color_data = 12'hfc5;
			{8'd102, 8'd32}: color_data = 12'h100;
			{8'd102, 8'd33}: color_data = 12'ha11;
			{8'd102, 8'd34}: color_data = 12'hf12;
			{8'd102, 8'd35}: color_data = 12'hf12;
			{8'd102, 8'd36}: color_data = 12'he12;
			{8'd102, 8'd37}: color_data = 12'he12;
			{8'd102, 8'd38}: color_data = 12'he12;
			{8'd102, 8'd39}: color_data = 12'he12;
			{8'd102, 8'd40}: color_data = 12'he12;
			{8'd102, 8'd41}: color_data = 12'he12;
			{8'd102, 8'd42}: color_data = 12'he12;
			{8'd102, 8'd43}: color_data = 12'he12;
			{8'd102, 8'd44}: color_data = 12'hf12;
			{8'd102, 8'd45}: color_data = 12'h934;
			{8'd102, 8'd46}: color_data = 12'hfff;
			{8'd102, 8'd47}: color_data = 12'hfff;
			{8'd102, 8'd48}: color_data = 12'hfbb;
			{8'd102, 8'd49}: color_data = 12'hfbc;
			{8'd102, 8'd50}: color_data = 12'heff;
			{8'd102, 8'd51}: color_data = 12'h934;
			{8'd102, 8'd52}: color_data = 12'hf11;
			{8'd102, 8'd53}: color_data = 12'he12;
			{8'd102, 8'd54}: color_data = 12'he12;
			{8'd102, 8'd55}: color_data = 12'h832;
			{8'd102, 8'd56}: color_data = 12'hcb9;
			{8'd102, 8'd57}: color_data = 12'hfdb;
			{8'd102, 8'd58}: color_data = 12'hfdb;
			{8'd102, 8'd59}: color_data = 12'hfda;
			{8'd102, 8'd60}: color_data = 12'hfda;
			{8'd102, 8'd61}: color_data = 12'hfdb;
			{8'd102, 8'd62}: color_data = 12'hfdb;
			{8'd102, 8'd63}: color_data = 12'hfdb;
			{8'd102, 8'd64}: color_data = 12'h986;
			{8'd102, 8'd65}: color_data = 12'h865;
			{8'd102, 8'd66}: color_data = 12'hfca;
			{8'd102, 8'd67}: color_data = 12'hfdb;
			{8'd102, 8'd68}: color_data = 12'hfdb;
			{8'd102, 8'd69}: color_data = 12'h865;
			{8'd102, 8'd70}: color_data = 12'h000;
			{8'd102, 8'd71}: color_data = 12'h000;
			{8'd102, 8'd72}: color_data = 12'h000;
			{8'd102, 8'd73}: color_data = 12'h000;
			{8'd102, 8'd74}: color_data = 12'h433;
			{8'd102, 8'd75}: color_data = 12'hfdb;
			{8'd102, 8'd76}: color_data = 12'hfdb;
			{8'd102, 8'd77}: color_data = 12'hfda;
			{8'd102, 8'd78}: color_data = 12'hfda;
			{8'd102, 8'd79}: color_data = 12'hfda;
			{8'd102, 8'd80}: color_data = 12'hfdb;
			{8'd102, 8'd81}: color_data = 12'ha87;
			{8'd102, 8'd82}: color_data = 12'h754;
			{8'd102, 8'd83}: color_data = 12'hccc;
			{8'd102, 8'd84}: color_data = 12'hfff;
			{8'd102, 8'd85}: color_data = 12'hfff;
			{8'd102, 8'd86}: color_data = 12'hfff;
			{8'd102, 8'd87}: color_data = 12'hfff;
			{8'd102, 8'd88}: color_data = 12'hfff;
			{8'd102, 8'd89}: color_data = 12'heee;
			{8'd102, 8'd90}: color_data = 12'hfff;
			{8'd102, 8'd91}: color_data = 12'hddd;
			{8'd102, 8'd92}: color_data = 12'hfff;
			{8'd102, 8'd93}: color_data = 12'hfff;
			{8'd102, 8'd94}: color_data = 12'hfff;
			{8'd102, 8'd95}: color_data = 12'hfff;
			{8'd102, 8'd96}: color_data = 12'hfff;
			{8'd102, 8'd97}: color_data = 12'hfff;
			{8'd102, 8'd98}: color_data = 12'h999;
			{8'd102, 8'd99}: color_data = 12'h755;
			{8'd102, 8'd100}: color_data = 12'hb86;
			{8'd102, 8'd101}: color_data = 12'hc97;
			{8'd102, 8'd102}: color_data = 12'hc97;
			{8'd102, 8'd103}: color_data = 12'hc97;
			{8'd102, 8'd104}: color_data = 12'h765;
			{8'd102, 8'd105}: color_data = 12'h047;
			{8'd102, 8'd106}: color_data = 12'h06b;
			{8'd102, 8'd107}: color_data = 12'h06b;
			{8'd102, 8'd108}: color_data = 12'h06b;
			{8'd102, 8'd109}: color_data = 12'h06b;
			{8'd102, 8'd110}: color_data = 12'h06b;
			{8'd102, 8'd111}: color_data = 12'h06b;
			{8'd102, 8'd112}: color_data = 12'h06b;
			{8'd102, 8'd113}: color_data = 12'h06b;
			{8'd102, 8'd114}: color_data = 12'h06b;
			{8'd102, 8'd115}: color_data = 12'h06b;
			{8'd102, 8'd116}: color_data = 12'h06b;
			{8'd102, 8'd117}: color_data = 12'h06b;
			{8'd102, 8'd118}: color_data = 12'h06b;
			{8'd102, 8'd119}: color_data = 12'h06b;
			{8'd102, 8'd120}: color_data = 12'h06b;
			{8'd102, 8'd121}: color_data = 12'h06b;
			{8'd102, 8'd122}: color_data = 12'h06b;
			{8'd102, 8'd123}: color_data = 12'h06b;
			{8'd102, 8'd124}: color_data = 12'h06b;
			{8'd102, 8'd125}: color_data = 12'h06b;
			{8'd102, 8'd126}: color_data = 12'h06b;
			{8'd102, 8'd127}: color_data = 12'h06b;
			{8'd102, 8'd128}: color_data = 12'h06b;
			{8'd102, 8'd129}: color_data = 12'h06b;
			{8'd102, 8'd130}: color_data = 12'h06b;
			{8'd102, 8'd131}: color_data = 12'h06b;
			{8'd102, 8'd132}: color_data = 12'h06b;
			{8'd102, 8'd133}: color_data = 12'h06b;
			{8'd102, 8'd134}: color_data = 12'h06b;
			{8'd102, 8'd135}: color_data = 12'h06b;
			{8'd102, 8'd136}: color_data = 12'h06b;
			{8'd102, 8'd137}: color_data = 12'h06b;
			{8'd102, 8'd138}: color_data = 12'h06b;
			{8'd102, 8'd139}: color_data = 12'h06b;
			{8'd102, 8'd140}: color_data = 12'h06b;
			{8'd102, 8'd141}: color_data = 12'h06b;
			{8'd102, 8'd142}: color_data = 12'h06b;
			{8'd102, 8'd143}: color_data = 12'h06b;
			{8'd102, 8'd144}: color_data = 12'h06b;
			{8'd102, 8'd145}: color_data = 12'h06b;
			{8'd102, 8'd146}: color_data = 12'h05a;
			{8'd102, 8'd147}: color_data = 12'h211;
			{8'd102, 8'd148}: color_data = 12'h842;
			{8'd102, 8'd149}: color_data = 12'h842;
			{8'd102, 8'd150}: color_data = 12'h842;
			{8'd102, 8'd151}: color_data = 12'h842;
			{8'd102, 8'd152}: color_data = 12'h842;
			{8'd102, 8'd153}: color_data = 12'h842;
			{8'd102, 8'd154}: color_data = 12'h842;
			{8'd102, 8'd155}: color_data = 12'h842;
			{8'd102, 8'd156}: color_data = 12'h842;
			{8'd102, 8'd157}: color_data = 12'h753;
			{8'd102, 8'd158}: color_data = 12'h532;
			{8'd103, 8'd3}: color_data = 12'hfc4;
			{8'd103, 8'd4}: color_data = 12'hfc5;
			{8'd103, 8'd5}: color_data = 12'hea1;
			{8'd103, 8'd6}: color_data = 12'hd90;
			{8'd103, 8'd7}: color_data = 12'hd90;
			{8'd103, 8'd8}: color_data = 12'hd90;
			{8'd103, 8'd9}: color_data = 12'hd90;
			{8'd103, 8'd10}: color_data = 12'hea2;
			{8'd103, 8'd11}: color_data = 12'heb3;
			{8'd103, 8'd12}: color_data = 12'hfb3;
			{8'd103, 8'd13}: color_data = 12'hea1;
			{8'd103, 8'd14}: color_data = 12'hd90;
			{8'd103, 8'd15}: color_data = 12'hd90;
			{8'd103, 8'd16}: color_data = 12'hd90;
			{8'd103, 8'd17}: color_data = 12'hd90;
			{8'd103, 8'd18}: color_data = 12'hd90;
			{8'd103, 8'd19}: color_data = 12'hfc4;
			{8'd103, 8'd20}: color_data = 12'hfc5;
			{8'd103, 8'd21}: color_data = 12'hfc5;
			{8'd103, 8'd33}: color_data = 12'h100;
			{8'd103, 8'd34}: color_data = 12'h701;
			{8'd103, 8'd35}: color_data = 12'hc11;
			{8'd103, 8'd36}: color_data = 12'he12;
			{8'd103, 8'd37}: color_data = 12'hf12;
			{8'd103, 8'd38}: color_data = 12'hf12;
			{8'd103, 8'd39}: color_data = 12'hf12;
			{8'd103, 8'd40}: color_data = 12'hf12;
			{8'd103, 8'd41}: color_data = 12'he12;
			{8'd103, 8'd42}: color_data = 12'he12;
			{8'd103, 8'd43}: color_data = 12'he12;
			{8'd103, 8'd44}: color_data = 12'hf12;
			{8'd103, 8'd45}: color_data = 12'hc12;
			{8'd103, 8'd46}: color_data = 12'ha88;
			{8'd103, 8'd47}: color_data = 12'hd88;
			{8'd103, 8'd48}: color_data = 12'hf88;
			{8'd103, 8'd49}: color_data = 12'hfdd;
			{8'd103, 8'd50}: color_data = 12'ha88;
			{8'd103, 8'd51}: color_data = 12'hc11;
			{8'd103, 8'd52}: color_data = 12'hf12;
			{8'd103, 8'd53}: color_data = 12'hf12;
			{8'd103, 8'd54}: color_data = 12'hb11;
			{8'd103, 8'd55}: color_data = 12'hc98;
			{8'd103, 8'd56}: color_data = 12'heca;
			{8'd103, 8'd57}: color_data = 12'hfca;
			{8'd103, 8'd58}: color_data = 12'hfdb;
			{8'd103, 8'd59}: color_data = 12'hfda;
			{8'd103, 8'd60}: color_data = 12'hfda;
			{8'd103, 8'd61}: color_data = 12'hfdb;
			{8'd103, 8'd62}: color_data = 12'hfca;
			{8'd103, 8'd63}: color_data = 12'h543;
			{8'd103, 8'd64}: color_data = 12'h322;
			{8'd103, 8'd65}: color_data = 12'hb97;
			{8'd103, 8'd66}: color_data = 12'hfca;
			{8'd103, 8'd67}: color_data = 12'hfda;
			{8'd103, 8'd68}: color_data = 12'hfdb;
			{8'd103, 8'd69}: color_data = 12'heca;
			{8'd103, 8'd70}: color_data = 12'h111;
			{8'd103, 8'd71}: color_data = 12'h000;
			{8'd103, 8'd72}: color_data = 12'h000;
			{8'd103, 8'd73}: color_data = 12'h000;
			{8'd103, 8'd74}: color_data = 12'h000;
			{8'd103, 8'd75}: color_data = 12'h755;
			{8'd103, 8'd76}: color_data = 12'hfca;
			{8'd103, 8'd77}: color_data = 12'hfdb;
			{8'd103, 8'd78}: color_data = 12'hfdb;
			{8'd103, 8'd79}: color_data = 12'hfdb;
			{8'd103, 8'd80}: color_data = 12'heba;
			{8'd103, 8'd81}: color_data = 12'h865;
			{8'd103, 8'd82}: color_data = 12'hc97;
			{8'd103, 8'd83}: color_data = 12'h865;
			{8'd103, 8'd84}: color_data = 12'haaa;
			{8'd103, 8'd85}: color_data = 12'hfff;
			{8'd103, 8'd86}: color_data = 12'hfff;
			{8'd103, 8'd87}: color_data = 12'hbbb;
			{8'd103, 8'd88}: color_data = 12'heee;
			{8'd103, 8'd89}: color_data = 12'hddd;
			{8'd103, 8'd90}: color_data = 12'haaa;
			{8'd103, 8'd91}: color_data = 12'hbbb;
			{8'd103, 8'd92}: color_data = 12'hddd;
			{8'd103, 8'd93}: color_data = 12'hfff;
			{8'd103, 8'd94}: color_data = 12'hfff;
			{8'd103, 8'd95}: color_data = 12'hfff;
			{8'd103, 8'd96}: color_data = 12'hfff;
			{8'd103, 8'd97}: color_data = 12'hfff;
			{8'd103, 8'd98}: color_data = 12'hbbb;
			{8'd103, 8'd99}: color_data = 12'hddd;
			{8'd103, 8'd100}: color_data = 12'h988;
			{8'd103, 8'd101}: color_data = 12'hb86;
			{8'd103, 8'd102}: color_data = 12'hc97;
			{8'd103, 8'd103}: color_data = 12'hc97;
			{8'd103, 8'd104}: color_data = 12'hd97;
			{8'd103, 8'd105}: color_data = 12'h965;
			{8'd103, 8'd106}: color_data = 12'h047;
			{8'd103, 8'd107}: color_data = 12'h06b;
			{8'd103, 8'd108}: color_data = 12'h06b;
			{8'd103, 8'd109}: color_data = 12'h06b;
			{8'd103, 8'd110}: color_data = 12'h06b;
			{8'd103, 8'd111}: color_data = 12'h06b;
			{8'd103, 8'd112}: color_data = 12'h06b;
			{8'd103, 8'd113}: color_data = 12'h06b;
			{8'd103, 8'd114}: color_data = 12'h06b;
			{8'd103, 8'd115}: color_data = 12'h05a;
			{8'd103, 8'd116}: color_data = 12'h059;
			{8'd103, 8'd117}: color_data = 12'h06b;
			{8'd103, 8'd118}: color_data = 12'h06b;
			{8'd103, 8'd119}: color_data = 12'h06b;
			{8'd103, 8'd120}: color_data = 12'h06b;
			{8'd103, 8'd121}: color_data = 12'h06b;
			{8'd103, 8'd122}: color_data = 12'h06b;
			{8'd103, 8'd123}: color_data = 12'h06b;
			{8'd103, 8'd124}: color_data = 12'h06b;
			{8'd103, 8'd125}: color_data = 12'h06b;
			{8'd103, 8'd126}: color_data = 12'h06b;
			{8'd103, 8'd127}: color_data = 12'h06b;
			{8'd103, 8'd128}: color_data = 12'h06b;
			{8'd103, 8'd129}: color_data = 12'h06b;
			{8'd103, 8'd130}: color_data = 12'h06b;
			{8'd103, 8'd131}: color_data = 12'h06b;
			{8'd103, 8'd132}: color_data = 12'h06b;
			{8'd103, 8'd133}: color_data = 12'h06b;
			{8'd103, 8'd134}: color_data = 12'h06b;
			{8'd103, 8'd135}: color_data = 12'h06b;
			{8'd103, 8'd136}: color_data = 12'h06b;
			{8'd103, 8'd137}: color_data = 12'h06b;
			{8'd103, 8'd138}: color_data = 12'h06b;
			{8'd103, 8'd139}: color_data = 12'h06b;
			{8'd103, 8'd140}: color_data = 12'h06b;
			{8'd103, 8'd141}: color_data = 12'h06b;
			{8'd103, 8'd142}: color_data = 12'h059;
			{8'd103, 8'd143}: color_data = 12'h035;
			{8'd103, 8'd144}: color_data = 12'h059;
			{8'd103, 8'd145}: color_data = 12'h05a;
			{8'd103, 8'd146}: color_data = 12'h036;
			{8'd103, 8'd147}: color_data = 12'h421;
			{8'd103, 8'd148}: color_data = 12'h843;
			{8'd103, 8'd149}: color_data = 12'h842;
			{8'd103, 8'd150}: color_data = 12'h842;
			{8'd103, 8'd151}: color_data = 12'h842;
			{8'd103, 8'd152}: color_data = 12'h842;
			{8'd103, 8'd153}: color_data = 12'h842;
			{8'd103, 8'd154}: color_data = 12'h842;
			{8'd103, 8'd155}: color_data = 12'h842;
			{8'd103, 8'd156}: color_data = 12'h842;
			{8'd103, 8'd157}: color_data = 12'h742;
			{8'd103, 8'd158}: color_data = 12'h542;
			{8'd104, 8'd2}: color_data = 12'hfc6;
			{8'd104, 8'd3}: color_data = 12'hfc4;
			{8'd104, 8'd4}: color_data = 12'hfc5;
			{8'd104, 8'd5}: color_data = 12'hea1;
			{8'd104, 8'd6}: color_data = 12'hd90;
			{8'd104, 8'd7}: color_data = 12'hd90;
			{8'd104, 8'd8}: color_data = 12'hd90;
			{8'd104, 8'd9}: color_data = 12'hfb3;
			{8'd104, 8'd10}: color_data = 12'hfd6;
			{8'd104, 8'd11}: color_data = 12'hfd6;
			{8'd104, 8'd12}: color_data = 12'hfd7;
			{8'd104, 8'd13}: color_data = 12'hfc6;
			{8'd104, 8'd14}: color_data = 12'heb2;
			{8'd104, 8'd15}: color_data = 12'hd90;
			{8'd104, 8'd16}: color_data = 12'hd90;
			{8'd104, 8'd17}: color_data = 12'hd90;
			{8'd104, 8'd18}: color_data = 12'hd90;
			{8'd104, 8'd19}: color_data = 12'hfc4;
			{8'd104, 8'd20}: color_data = 12'hfc5;
			{8'd104, 8'd21}: color_data = 12'hfc6;
			{8'd104, 8'd34}: color_data = 12'h000;
			{8'd104, 8'd35}: color_data = 12'h100;
			{8'd104, 8'd36}: color_data = 12'h500;
			{8'd104, 8'd37}: color_data = 12'h801;
			{8'd104, 8'd38}: color_data = 12'ha11;
			{8'd104, 8'd39}: color_data = 12'hc11;
			{8'd104, 8'd40}: color_data = 12'hd12;
			{8'd104, 8'd41}: color_data = 12'he12;
			{8'd104, 8'd42}: color_data = 12'hf12;
			{8'd104, 8'd43}: color_data = 12'hf12;
			{8'd104, 8'd44}: color_data = 12'hf12;
			{8'd104, 8'd45}: color_data = 12'hf12;
			{8'd104, 8'd46}: color_data = 12'hd11;
			{8'd104, 8'd47}: color_data = 12'ha22;
			{8'd104, 8'd48}: color_data = 12'h833;
			{8'd104, 8'd49}: color_data = 12'h633;
			{8'd104, 8'd50}: color_data = 12'h811;
			{8'd104, 8'd51}: color_data = 12'hf12;
			{8'd104, 8'd52}: color_data = 12'he12;
			{8'd104, 8'd53}: color_data = 12'he12;
			{8'd104, 8'd54}: color_data = 12'h632;
			{8'd104, 8'd55}: color_data = 12'hfdb;
			{8'd104, 8'd56}: color_data = 12'hca8;
			{8'd104, 8'd57}: color_data = 12'h986;
			{8'd104, 8'd58}: color_data = 12'heb9;
			{8'd104, 8'd59}: color_data = 12'hfdb;
			{8'd104, 8'd60}: color_data = 12'hfdb;
			{8'd104, 8'd61}: color_data = 12'hfca;
			{8'd104, 8'd62}: color_data = 12'h433;
			{8'd104, 8'd63}: color_data = 12'h433;
			{8'd104, 8'd64}: color_data = 12'hfca;
			{8'd104, 8'd65}: color_data = 12'hfdb;
			{8'd104, 8'd66}: color_data = 12'hfda;
			{8'd104, 8'd67}: color_data = 12'hfda;
			{8'd104, 8'd68}: color_data = 12'hfda;
			{8'd104, 8'd69}: color_data = 12'hfdb;
			{8'd104, 8'd70}: color_data = 12'h765;
			{8'd104, 8'd71}: color_data = 12'h000;
			{8'd104, 8'd72}: color_data = 12'h000;
			{8'd104, 8'd73}: color_data = 12'h000;
			{8'd104, 8'd74}: color_data = 12'h000;
			{8'd104, 8'd75}: color_data = 12'h000;
			{8'd104, 8'd76}: color_data = 12'ha87;
			{8'd104, 8'd77}: color_data = 12'hfdb;
			{8'd104, 8'd78}: color_data = 12'hfca;
			{8'd104, 8'd79}: color_data = 12'hfdb;
			{8'd104, 8'd80}: color_data = 12'h765;
			{8'd104, 8'd81}: color_data = 12'ha86;
			{8'd104, 8'd82}: color_data = 12'hc97;
			{8'd104, 8'd83}: color_data = 12'hc97;
			{8'd104, 8'd84}: color_data = 12'ha76;
			{8'd104, 8'd85}: color_data = 12'h877;
			{8'd104, 8'd86}: color_data = 12'hbbb;
			{8'd104, 8'd87}: color_data = 12'hddd;
			{8'd104, 8'd88}: color_data = 12'haaa;
			{8'd104, 8'd89}: color_data = 12'hfff;
			{8'd104, 8'd90}: color_data = 12'hccc;
			{8'd104, 8'd91}: color_data = 12'heee;
			{8'd104, 8'd92}: color_data = 12'hfff;
			{8'd104, 8'd93}: color_data = 12'hfff;
			{8'd104, 8'd94}: color_data = 12'hfff;
			{8'd104, 8'd95}: color_data = 12'hfff;
			{8'd104, 8'd96}: color_data = 12'hfff;
			{8'd104, 8'd97}: color_data = 12'hfff;
			{8'd104, 8'd98}: color_data = 12'haaa;
			{8'd104, 8'd99}: color_data = 12'hfff;
			{8'd104, 8'd100}: color_data = 12'hddd;
			{8'd104, 8'd101}: color_data = 12'h975;
			{8'd104, 8'd102}: color_data = 12'hc97;
			{8'd104, 8'd103}: color_data = 12'hc97;
			{8'd104, 8'd104}: color_data = 12'hc97;
			{8'd104, 8'd105}: color_data = 12'hd97;
			{8'd104, 8'd106}: color_data = 12'h865;
			{8'd104, 8'd107}: color_data = 12'h048;
			{8'd104, 8'd108}: color_data = 12'h06b;
			{8'd104, 8'd109}: color_data = 12'h06b;
			{8'd104, 8'd110}: color_data = 12'h06b;
			{8'd104, 8'd111}: color_data = 12'h06b;
			{8'd104, 8'd112}: color_data = 12'h06b;
			{8'd104, 8'd113}: color_data = 12'h05a;
			{8'd104, 8'd114}: color_data = 12'h048;
			{8'd104, 8'd115}: color_data = 12'h555;
			{8'd104, 8'd116}: color_data = 12'h765;
			{8'd104, 8'd117}: color_data = 12'h246;
			{8'd104, 8'd118}: color_data = 12'h059;
			{8'd104, 8'd119}: color_data = 12'h06b;
			{8'd104, 8'd120}: color_data = 12'h06b;
			{8'd104, 8'd121}: color_data = 12'h06b;
			{8'd104, 8'd122}: color_data = 12'h06b;
			{8'd104, 8'd123}: color_data = 12'h06b;
			{8'd104, 8'd124}: color_data = 12'h06b;
			{8'd104, 8'd125}: color_data = 12'h06b;
			{8'd104, 8'd126}: color_data = 12'h06b;
			{8'd104, 8'd127}: color_data = 12'h06b;
			{8'd104, 8'd128}: color_data = 12'h06b;
			{8'd104, 8'd129}: color_data = 12'h06b;
			{8'd104, 8'd130}: color_data = 12'h06b;
			{8'd104, 8'd131}: color_data = 12'h06b;
			{8'd104, 8'd132}: color_data = 12'h06b;
			{8'd104, 8'd133}: color_data = 12'h06b;
			{8'd104, 8'd134}: color_data = 12'h06b;
			{8'd104, 8'd135}: color_data = 12'h06b;
			{8'd104, 8'd136}: color_data = 12'h06b;
			{8'd104, 8'd137}: color_data = 12'h06b;
			{8'd104, 8'd138}: color_data = 12'h06b;
			{8'd104, 8'd139}: color_data = 12'h06b;
			{8'd104, 8'd140}: color_data = 12'h06b;
			{8'd104, 8'd141}: color_data = 12'h06a;
			{8'd104, 8'd142}: color_data = 12'h023;
			{8'd104, 8'd143}: color_data = 12'h000;
			{8'd104, 8'd144}: color_data = 12'h012;
			{8'd104, 8'd145}: color_data = 12'h012;
			{8'd104, 8'd146}: color_data = 12'h000;
			{8'd104, 8'd147}: color_data = 12'h521;
			{8'd104, 8'd148}: color_data = 12'h843;
			{8'd104, 8'd149}: color_data = 12'h842;
			{8'd104, 8'd150}: color_data = 12'h842;
			{8'd104, 8'd151}: color_data = 12'h842;
			{8'd104, 8'd152}: color_data = 12'h842;
			{8'd104, 8'd153}: color_data = 12'h842;
			{8'd104, 8'd154}: color_data = 12'h842;
			{8'd104, 8'd155}: color_data = 12'h842;
			{8'd104, 8'd156}: color_data = 12'h843;
			{8'd104, 8'd157}: color_data = 12'h742;
			{8'd104, 8'd158}: color_data = 12'h542;
			{8'd105, 8'd2}: color_data = 12'hec5;
			{8'd105, 8'd3}: color_data = 12'hfc5;
			{8'd105, 8'd4}: color_data = 12'hfc4;
			{8'd105, 8'd5}: color_data = 12'hea0;
			{8'd105, 8'd6}: color_data = 12'hd90;
			{8'd105, 8'd7}: color_data = 12'hd90;
			{8'd105, 8'd8}: color_data = 12'hea0;
			{8'd105, 8'd9}: color_data = 12'hfc5;
			{8'd105, 8'd10}: color_data = 12'heb2;
			{8'd105, 8'd11}: color_data = 12'hea1;
			{8'd105, 8'd12}: color_data = 12'heb2;
			{8'd105, 8'd13}: color_data = 12'hfb4;
			{8'd105, 8'd14}: color_data = 12'hfc4;
			{8'd105, 8'd15}: color_data = 12'hd90;
			{8'd105, 8'd16}: color_data = 12'hd90;
			{8'd105, 8'd17}: color_data = 12'hd90;
			{8'd105, 8'd18}: color_data = 12'hea1;
			{8'd105, 8'd19}: color_data = 12'hfc5;
			{8'd105, 8'd20}: color_data = 12'hfc5;
			{8'd105, 8'd21}: color_data = 12'hff7;
			{8'd105, 8'd37}: color_data = 12'h000;
			{8'd105, 8'd38}: color_data = 12'h000;
			{8'd105, 8'd39}: color_data = 12'h100;
			{8'd105, 8'd40}: color_data = 12'h300;
			{8'd105, 8'd41}: color_data = 12'h400;
			{8'd105, 8'd42}: color_data = 12'h500;
			{8'd105, 8'd43}: color_data = 12'h600;
			{8'd105, 8'd44}: color_data = 12'h601;
			{8'd105, 8'd45}: color_data = 12'h600;
			{8'd105, 8'd46}: color_data = 12'h600;
			{8'd105, 8'd47}: color_data = 12'h500;
			{8'd105, 8'd48}: color_data = 12'h300;
			{8'd105, 8'd49}: color_data = 12'h200;
			{8'd105, 8'd50}: color_data = 12'hd11;
			{8'd105, 8'd51}: color_data = 12'hf12;
			{8'd105, 8'd52}: color_data = 12'hf12;
			{8'd105, 8'd53}: color_data = 12'ha11;
			{8'd105, 8'd54}: color_data = 12'h000;
			{8'd105, 8'd55}: color_data = 12'h765;
			{8'd105, 8'd56}: color_data = 12'hfca;
			{8'd105, 8'd57}: color_data = 12'heca;
			{8'd105, 8'd58}: color_data = 12'ha87;
			{8'd105, 8'd59}: color_data = 12'h986;
			{8'd105, 8'd60}: color_data = 12'hb98;
			{8'd105, 8'd61}: color_data = 12'hda9;
			{8'd105, 8'd62}: color_data = 12'h211;
			{8'd105, 8'd63}: color_data = 12'heb9;
			{8'd105, 8'd64}: color_data = 12'hfdb;
			{8'd105, 8'd65}: color_data = 12'hfda;
			{8'd105, 8'd66}: color_data = 12'hfda;
			{8'd105, 8'd67}: color_data = 12'hfda;
			{8'd105, 8'd68}: color_data = 12'hfda;
			{8'd105, 8'd69}: color_data = 12'hfdb;
			{8'd105, 8'd70}: color_data = 12'hb98;
			{8'd105, 8'd71}: color_data = 12'h000;
			{8'd105, 8'd72}: color_data = 12'h000;
			{8'd105, 8'd73}: color_data = 12'h000;
			{8'd105, 8'd74}: color_data = 12'h000;
			{8'd105, 8'd75}: color_data = 12'h000;
			{8'd105, 8'd76}: color_data = 12'h976;
			{8'd105, 8'd77}: color_data = 12'hca8;
			{8'd105, 8'd78}: color_data = 12'hdb9;
			{8'd105, 8'd79}: color_data = 12'h987;
			{8'd105, 8'd80}: color_data = 12'h112;
			{8'd105, 8'd81}: color_data = 12'ha76;
			{8'd105, 8'd82}: color_data = 12'hc97;
			{8'd105, 8'd83}: color_data = 12'hc97;
			{8'd105, 8'd84}: color_data = 12'hc97;
			{8'd105, 8'd85}: color_data = 12'h843;
			{8'd105, 8'd86}: color_data = 12'h801;
			{8'd105, 8'd87}: color_data = 12'h999;
			{8'd105, 8'd88}: color_data = 12'haaa;
			{8'd105, 8'd89}: color_data = 12'h777;
			{8'd105, 8'd90}: color_data = 12'h999;
			{8'd105, 8'd91}: color_data = 12'hddd;
			{8'd105, 8'd92}: color_data = 12'hfff;
			{8'd105, 8'd93}: color_data = 12'hfff;
			{8'd105, 8'd94}: color_data = 12'heee;
			{8'd105, 8'd95}: color_data = 12'hfff;
			{8'd105, 8'd96}: color_data = 12'hfff;
			{8'd105, 8'd97}: color_data = 12'hfff;
			{8'd105, 8'd98}: color_data = 12'hfff;
			{8'd105, 8'd99}: color_data = 12'hfff;
			{8'd105, 8'd100}: color_data = 12'h999;
			{8'd105, 8'd101}: color_data = 12'h643;
			{8'd105, 8'd102}: color_data = 12'hb86;
			{8'd105, 8'd103}: color_data = 12'hc97;
			{8'd105, 8'd104}: color_data = 12'hc97;
			{8'd105, 8'd105}: color_data = 12'hc97;
			{8'd105, 8'd106}: color_data = 12'hd97;
			{8'd105, 8'd107}: color_data = 12'h555;
			{8'd105, 8'd108}: color_data = 12'h048;
			{8'd105, 8'd109}: color_data = 12'h048;
			{8'd105, 8'd110}: color_data = 12'h047;
			{8'd105, 8'd111}: color_data = 12'h147;
			{8'd105, 8'd112}: color_data = 12'h346;
			{8'd105, 8'd113}: color_data = 12'h655;
			{8'd105, 8'd114}: color_data = 12'ha76;
			{8'd105, 8'd115}: color_data = 12'hc97;
			{8'd105, 8'd116}: color_data = 12'hd97;
			{8'd105, 8'd117}: color_data = 12'hc86;
			{8'd105, 8'd118}: color_data = 12'h765;
			{8'd105, 8'd119}: color_data = 12'h246;
			{8'd105, 8'd120}: color_data = 12'h058;
			{8'd105, 8'd121}: color_data = 12'h06a;
			{8'd105, 8'd122}: color_data = 12'h06b;
			{8'd105, 8'd123}: color_data = 12'h06b;
			{8'd105, 8'd124}: color_data = 12'h06b;
			{8'd105, 8'd125}: color_data = 12'h06b;
			{8'd105, 8'd126}: color_data = 12'h06b;
			{8'd105, 8'd127}: color_data = 12'h06b;
			{8'd105, 8'd128}: color_data = 12'h06b;
			{8'd105, 8'd129}: color_data = 12'h06b;
			{8'd105, 8'd130}: color_data = 12'h06b;
			{8'd105, 8'd131}: color_data = 12'h06b;
			{8'd105, 8'd132}: color_data = 12'h06b;
			{8'd105, 8'd133}: color_data = 12'h06b;
			{8'd105, 8'd134}: color_data = 12'h06b;
			{8'd105, 8'd135}: color_data = 12'h06b;
			{8'd105, 8'd136}: color_data = 12'h06b;
			{8'd105, 8'd137}: color_data = 12'h06b;
			{8'd105, 8'd138}: color_data = 12'h06b;
			{8'd105, 8'd139}: color_data = 12'h06b;
			{8'd105, 8'd140}: color_data = 12'h06b;
			{8'd105, 8'd141}: color_data = 12'h025;
			{8'd105, 8'd142}: color_data = 12'h000;
			{8'd105, 8'd147}: color_data = 12'h421;
			{8'd105, 8'd148}: color_data = 12'h843;
			{8'd105, 8'd149}: color_data = 12'h842;
			{8'd105, 8'd150}: color_data = 12'h842;
			{8'd105, 8'd151}: color_data = 12'h842;
			{8'd105, 8'd152}: color_data = 12'h842;
			{8'd105, 8'd153}: color_data = 12'h842;
			{8'd105, 8'd154}: color_data = 12'h842;
			{8'd105, 8'd155}: color_data = 12'h842;
			{8'd105, 8'd156}: color_data = 12'h843;
			{8'd105, 8'd157}: color_data = 12'h742;
			{8'd105, 8'd158}: color_data = 12'h542;
			{8'd105, 8'd159}: color_data = 12'h000;
			{8'd106, 8'd2}: color_data = 12'hfc5;
			{8'd106, 8'd3}: color_data = 12'hfc5;
			{8'd106, 8'd4}: color_data = 12'hfc4;
			{8'd106, 8'd5}: color_data = 12'hd90;
			{8'd106, 8'd6}: color_data = 12'hd90;
			{8'd106, 8'd7}: color_data = 12'hd90;
			{8'd106, 8'd8}: color_data = 12'hd90;
			{8'd106, 8'd9}: color_data = 12'hfc4;
			{8'd106, 8'd10}: color_data = 12'hda0;
			{8'd106, 8'd11}: color_data = 12'hd90;
			{8'd106, 8'd12}: color_data = 12'hd90;
			{8'd106, 8'd13}: color_data = 12'heb2;
			{8'd106, 8'd14}: color_data = 12'heb2;
			{8'd106, 8'd15}: color_data = 12'hd90;
			{8'd106, 8'd16}: color_data = 12'hd90;
			{8'd106, 8'd17}: color_data = 12'hd90;
			{8'd106, 8'd18}: color_data = 12'hfb3;
			{8'd106, 8'd19}: color_data = 12'hfc5;
			{8'd106, 8'd20}: color_data = 12'hfc5;
			{8'd106, 8'd48}: color_data = 12'h000;
			{8'd106, 8'd49}: color_data = 12'h811;
			{8'd106, 8'd50}: color_data = 12'hf12;
			{8'd106, 8'd51}: color_data = 12'hf12;
			{8'd106, 8'd52}: color_data = 12'hd12;
			{8'd106, 8'd53}: color_data = 12'h300;
			{8'd106, 8'd55}: color_data = 12'h000;
			{8'd106, 8'd56}: color_data = 12'h543;
			{8'd106, 8'd57}: color_data = 12'hca8;
			{8'd106, 8'd58}: color_data = 12'hfdb;
			{8'd106, 8'd59}: color_data = 12'hfca;
			{8'd106, 8'd60}: color_data = 12'heca;
			{8'd106, 8'd61}: color_data = 12'hfca;
			{8'd106, 8'd62}: color_data = 12'hca8;
			{8'd106, 8'd63}: color_data = 12'hfda;
			{8'd106, 8'd64}: color_data = 12'hfda;
			{8'd106, 8'd65}: color_data = 12'hfda;
			{8'd106, 8'd66}: color_data = 12'hfda;
			{8'd106, 8'd67}: color_data = 12'hfda;
			{8'd106, 8'd68}: color_data = 12'hfda;
			{8'd106, 8'd69}: color_data = 12'hfdb;
			{8'd106, 8'd70}: color_data = 12'hca8;
			{8'd106, 8'd71}: color_data = 12'h000;
			{8'd106, 8'd72}: color_data = 12'h000;
			{8'd106, 8'd73}: color_data = 12'h000;
			{8'd106, 8'd74}: color_data = 12'h000;
			{8'd106, 8'd75}: color_data = 12'h000;
			{8'd106, 8'd76}: color_data = 12'ha87;
			{8'd106, 8'd77}: color_data = 12'ha97;
			{8'd106, 8'd78}: color_data = 12'h654;
			{8'd106, 8'd79}: color_data = 12'h123;
			{8'd106, 8'd80}: color_data = 12'h124;
			{8'd106, 8'd81}: color_data = 12'h865;
			{8'd106, 8'd82}: color_data = 12'hc97;
			{8'd106, 8'd83}: color_data = 12'hc97;
			{8'd106, 8'd84}: color_data = 12'h975;
			{8'd106, 8'd85}: color_data = 12'hb11;
			{8'd106, 8'd86}: color_data = 12'hc12;
			{8'd106, 8'd87}: color_data = 12'hcdd;
			{8'd106, 8'd88}: color_data = 12'hfff;
			{8'd106, 8'd89}: color_data = 12'hccc;
			{8'd106, 8'd90}: color_data = 12'h999;
			{8'd106, 8'd91}: color_data = 12'h999;
			{8'd106, 8'd92}: color_data = 12'haaa;
			{8'd106, 8'd93}: color_data = 12'haaa;
			{8'd106, 8'd94}: color_data = 12'haaa;
			{8'd106, 8'd95}: color_data = 12'heee;
			{8'd106, 8'd96}: color_data = 12'hfff;
			{8'd106, 8'd97}: color_data = 12'hfff;
			{8'd106, 8'd98}: color_data = 12'hfff;
			{8'd106, 8'd99}: color_data = 12'haaa;
			{8'd106, 8'd100}: color_data = 12'h975;
			{8'd106, 8'd101}: color_data = 12'hb97;
			{8'd106, 8'd102}: color_data = 12'h754;
			{8'd106, 8'd103}: color_data = 12'hb86;
			{8'd106, 8'd104}: color_data = 12'hc97;
			{8'd106, 8'd105}: color_data = 12'hc97;
			{8'd106, 8'd106}: color_data = 12'hc97;
			{8'd106, 8'd107}: color_data = 12'hb86;
			{8'd106, 8'd108}: color_data = 12'h643;
			{8'd106, 8'd109}: color_data = 12'ha76;
			{8'd106, 8'd110}: color_data = 12'hb86;
			{8'd106, 8'd111}: color_data = 12'hb86;
			{8'd106, 8'd112}: color_data = 12'hc97;
			{8'd106, 8'd113}: color_data = 12'hd97;
			{8'd106, 8'd114}: color_data = 12'hc97;
			{8'd106, 8'd115}: color_data = 12'hc97;
			{8'd106, 8'd116}: color_data = 12'hc97;
			{8'd106, 8'd117}: color_data = 12'hc97;
			{8'd106, 8'd118}: color_data = 12'hd97;
			{8'd106, 8'd119}: color_data = 12'hc97;
			{8'd106, 8'd120}: color_data = 12'h975;
			{8'd106, 8'd121}: color_data = 12'h455;
			{8'd106, 8'd122}: color_data = 12'h147;
			{8'd106, 8'd123}: color_data = 12'h059;
			{8'd106, 8'd124}: color_data = 12'h06b;
			{8'd106, 8'd125}: color_data = 12'h06b;
			{8'd106, 8'd126}: color_data = 12'h06b;
			{8'd106, 8'd127}: color_data = 12'h06b;
			{8'd106, 8'd128}: color_data = 12'h06b;
			{8'd106, 8'd129}: color_data = 12'h06b;
			{8'd106, 8'd130}: color_data = 12'h06b;
			{8'd106, 8'd131}: color_data = 12'h06b;
			{8'd106, 8'd132}: color_data = 12'h06b;
			{8'd106, 8'd133}: color_data = 12'h06b;
			{8'd106, 8'd134}: color_data = 12'h06b;
			{8'd106, 8'd135}: color_data = 12'h06b;
			{8'd106, 8'd136}: color_data = 12'h06b;
			{8'd106, 8'd137}: color_data = 12'h06b;
			{8'd106, 8'd138}: color_data = 12'h06b;
			{8'd106, 8'd139}: color_data = 12'h06a;
			{8'd106, 8'd140}: color_data = 12'h025;
			{8'd106, 8'd141}: color_data = 12'h000;
			{8'd106, 8'd147}: color_data = 12'h311;
			{8'd106, 8'd148}: color_data = 12'h842;
			{8'd106, 8'd149}: color_data = 12'h842;
			{8'd106, 8'd150}: color_data = 12'h842;
			{8'd106, 8'd151}: color_data = 12'h842;
			{8'd106, 8'd152}: color_data = 12'h842;
			{8'd106, 8'd153}: color_data = 12'h842;
			{8'd106, 8'd154}: color_data = 12'h842;
			{8'd106, 8'd155}: color_data = 12'h842;
			{8'd106, 8'd156}: color_data = 12'h843;
			{8'd106, 8'd157}: color_data = 12'h742;
			{8'd106, 8'd158}: color_data = 12'h542;
			{8'd106, 8'd159}: color_data = 12'h000;
			{8'd107, 8'd2}: color_data = 12'heb4;
			{8'd107, 8'd3}: color_data = 12'hfc5;
			{8'd107, 8'd4}: color_data = 12'hfc5;
			{8'd107, 8'd5}: color_data = 12'hda0;
			{8'd107, 8'd6}: color_data = 12'hd90;
			{8'd107, 8'd7}: color_data = 12'hd90;
			{8'd107, 8'd8}: color_data = 12'hea1;
			{8'd107, 8'd9}: color_data = 12'hfb3;
			{8'd107, 8'd10}: color_data = 12'hd90;
			{8'd107, 8'd11}: color_data = 12'hd90;
			{8'd107, 8'd12}: color_data = 12'hd90;
			{8'd107, 8'd13}: color_data = 12'hfb2;
			{8'd107, 8'd14}: color_data = 12'hda0;
			{8'd107, 8'd15}: color_data = 12'hd90;
			{8'd107, 8'd16}: color_data = 12'hd90;
			{8'd107, 8'd17}: color_data = 12'hda0;
			{8'd107, 8'd18}: color_data = 12'hfc5;
			{8'd107, 8'd19}: color_data = 12'hfc5;
			{8'd107, 8'd20}: color_data = 12'hfc5;
			{8'd107, 8'd48}: color_data = 12'h300;
			{8'd107, 8'd49}: color_data = 12'hd12;
			{8'd107, 8'd50}: color_data = 12'hf12;
			{8'd107, 8'd51}: color_data = 12'hf12;
			{8'd107, 8'd52}: color_data = 12'h701;
			{8'd107, 8'd53}: color_data = 12'h000;
			{8'd107, 8'd56}: color_data = 12'h000;
			{8'd107, 8'd57}: color_data = 12'h000;
			{8'd107, 8'd58}: color_data = 12'h654;
			{8'd107, 8'd59}: color_data = 12'hda9;
			{8'd107, 8'd60}: color_data = 12'hfca;
			{8'd107, 8'd61}: color_data = 12'hfdb;
			{8'd107, 8'd62}: color_data = 12'hfca;
			{8'd107, 8'd63}: color_data = 12'hca8;
			{8'd107, 8'd64}: color_data = 12'hfda;
			{8'd107, 8'd65}: color_data = 12'hfda;
			{8'd107, 8'd66}: color_data = 12'hfda;
			{8'd107, 8'd67}: color_data = 12'hfda;
			{8'd107, 8'd68}: color_data = 12'hfda;
			{8'd107, 8'd69}: color_data = 12'hfdb;
			{8'd107, 8'd70}: color_data = 12'h765;
			{8'd107, 8'd71}: color_data = 12'h000;
			{8'd107, 8'd72}: color_data = 12'h000;
			{8'd107, 8'd73}: color_data = 12'h000;
			{8'd107, 8'd74}: color_data = 12'h000;
			{8'd107, 8'd75}: color_data = 12'h100;
			{8'd107, 8'd76}: color_data = 12'heb9;
			{8'd107, 8'd77}: color_data = 12'h976;
			{8'd107, 8'd78}: color_data = 12'h754;
			{8'd107, 8'd79}: color_data = 12'h123;
			{8'd107, 8'd80}: color_data = 12'h134;
			{8'd107, 8'd81}: color_data = 12'h544;
			{8'd107, 8'd82}: color_data = 12'hc97;
			{8'd107, 8'd83}: color_data = 12'hc97;
			{8'd107, 8'd84}: color_data = 12'h832;
			{8'd107, 8'd85}: color_data = 12'hf12;
			{8'd107, 8'd86}: color_data = 12'hd11;
			{8'd107, 8'd87}: color_data = 12'h977;
			{8'd107, 8'd88}: color_data = 12'hfff;
			{8'd107, 8'd89}: color_data = 12'hfff;
			{8'd107, 8'd90}: color_data = 12'hfff;
			{8'd107, 8'd91}: color_data = 12'hfff;
			{8'd107, 8'd92}: color_data = 12'hfff;
			{8'd107, 8'd93}: color_data = 12'hfff;
			{8'd107, 8'd94}: color_data = 12'hfff;
			{8'd107, 8'd95}: color_data = 12'hfff;
			{8'd107, 8'd96}: color_data = 12'hfff;
			{8'd107, 8'd97}: color_data = 12'heee;
			{8'd107, 8'd98}: color_data = 12'ha88;
			{8'd107, 8'd99}: color_data = 12'h811;
			{8'd107, 8'd100}: color_data = 12'ha75;
			{8'd107, 8'd101}: color_data = 12'hd97;
			{8'd107, 8'd102}: color_data = 12'hc97;
			{8'd107, 8'd103}: color_data = 12'h754;
			{8'd107, 8'd104}: color_data = 12'hb87;
			{8'd107, 8'd105}: color_data = 12'hc97;
			{8'd107, 8'd106}: color_data = 12'hc97;
			{8'd107, 8'd107}: color_data = 12'hc97;
			{8'd107, 8'd108}: color_data = 12'ha86;
			{8'd107, 8'd109}: color_data = 12'hc97;
			{8'd107, 8'd110}: color_data = 12'hc97;
			{8'd107, 8'd111}: color_data = 12'hc97;
			{8'd107, 8'd112}: color_data = 12'hc97;
			{8'd107, 8'd113}: color_data = 12'hc97;
			{8'd107, 8'd114}: color_data = 12'hc97;
			{8'd107, 8'd115}: color_data = 12'hc97;
			{8'd107, 8'd116}: color_data = 12'hc97;
			{8'd107, 8'd117}: color_data = 12'hc97;
			{8'd107, 8'd118}: color_data = 12'hc97;
			{8'd107, 8'd119}: color_data = 12'hc97;
			{8'd107, 8'd120}: color_data = 12'hc97;
			{8'd107, 8'd121}: color_data = 12'hc97;
			{8'd107, 8'd122}: color_data = 12'hb86;
			{8'd107, 8'd123}: color_data = 12'h865;
			{8'd107, 8'd124}: color_data = 12'h455;
			{8'd107, 8'd125}: color_data = 12'h147;
			{8'd107, 8'd126}: color_data = 12'h058;
			{8'd107, 8'd127}: color_data = 12'h05a;
			{8'd107, 8'd128}: color_data = 12'h06b;
			{8'd107, 8'd129}: color_data = 12'h06b;
			{8'd107, 8'd130}: color_data = 12'h06b;
			{8'd107, 8'd131}: color_data = 12'h06b;
			{8'd107, 8'd132}: color_data = 12'h06b;
			{8'd107, 8'd133}: color_data = 12'h06b;
			{8'd107, 8'd134}: color_data = 12'h06b;
			{8'd107, 8'd135}: color_data = 12'h06b;
			{8'd107, 8'd136}: color_data = 12'h06b;
			{8'd107, 8'd137}: color_data = 12'h06b;
			{8'd107, 8'd138}: color_data = 12'h059;
			{8'd107, 8'd139}: color_data = 12'h024;
			{8'd107, 8'd140}: color_data = 12'h000;
			{8'd107, 8'd147}: color_data = 12'h100;
			{8'd107, 8'd148}: color_data = 12'h742;
			{8'd107, 8'd149}: color_data = 12'h843;
			{8'd107, 8'd150}: color_data = 12'h842;
			{8'd107, 8'd151}: color_data = 12'h842;
			{8'd107, 8'd152}: color_data = 12'h842;
			{8'd107, 8'd153}: color_data = 12'h842;
			{8'd107, 8'd154}: color_data = 12'h842;
			{8'd107, 8'd155}: color_data = 12'h842;
			{8'd107, 8'd156}: color_data = 12'h842;
			{8'd107, 8'd157}: color_data = 12'h742;
			{8'd107, 8'd158}: color_data = 12'h642;
			{8'd108, 8'd2}: color_data = 12'hfb4;
			{8'd108, 8'd3}: color_data = 12'hfc4;
			{8'd108, 8'd4}: color_data = 12'hfc5;
			{8'd108, 8'd5}: color_data = 12'hfb3;
			{8'd108, 8'd6}: color_data = 12'hd90;
			{8'd108, 8'd7}: color_data = 12'hea0;
			{8'd108, 8'd8}: color_data = 12'hfc6;
			{8'd108, 8'd9}: color_data = 12'heb3;
			{8'd108, 8'd10}: color_data = 12'hd90;
			{8'd108, 8'd11}: color_data = 12'hd90;
			{8'd108, 8'd12}: color_data = 12'hd90;
			{8'd108, 8'd13}: color_data = 12'hda0;
			{8'd108, 8'd14}: color_data = 12'hd90;
			{8'd108, 8'd15}: color_data = 12'hd90;
			{8'd108, 8'd16}: color_data = 12'hd90;
			{8'd108, 8'd17}: color_data = 12'hea1;
			{8'd108, 8'd18}: color_data = 12'hfc5;
			{8'd108, 8'd19}: color_data = 12'hfc5;
			{8'd108, 8'd47}: color_data = 12'h000;
			{8'd108, 8'd48}: color_data = 12'h911;
			{8'd108, 8'd49}: color_data = 12'hf12;
			{8'd108, 8'd50}: color_data = 12'hf12;
			{8'd108, 8'd51}: color_data = 12'ha11;
			{8'd108, 8'd52}: color_data = 12'h000;
			{8'd108, 8'd54}: color_data = 12'h000;
			{8'd108, 8'd55}: color_data = 12'h321;
			{8'd108, 8'd56}: color_data = 12'hb94;
			{8'd108, 8'd57}: color_data = 12'ha84;
			{8'd108, 8'd58}: color_data = 12'ha94;
			{8'd108, 8'd59}: color_data = 12'h974;
			{8'd108, 8'd60}: color_data = 12'h975;
			{8'd108, 8'd61}: color_data = 12'ha86;
			{8'd108, 8'd62}: color_data = 12'h976;
			{8'd108, 8'd63}: color_data = 12'hdb9;
			{8'd108, 8'd64}: color_data = 12'hfdb;
			{8'd108, 8'd65}: color_data = 12'hfda;
			{8'd108, 8'd66}: color_data = 12'hfda;
			{8'd108, 8'd67}: color_data = 12'hfda;
			{8'd108, 8'd68}: color_data = 12'hfda;
			{8'd108, 8'd69}: color_data = 12'hfdb;
			{8'd108, 8'd70}: color_data = 12'hca8;
			{8'd108, 8'd71}: color_data = 12'h000;
			{8'd108, 8'd72}: color_data = 12'h000;
			{8'd108, 8'd73}: color_data = 12'h000;
			{8'd108, 8'd74}: color_data = 12'h000;
			{8'd108, 8'd75}: color_data = 12'h221;
			{8'd108, 8'd76}: color_data = 12'heca;
			{8'd108, 8'd77}: color_data = 12'h975;
			{8'd108, 8'd78}: color_data = 12'h765;
			{8'd108, 8'd79}: color_data = 12'h113;
			{8'd108, 8'd80}: color_data = 12'h124;
			{8'd108, 8'd81}: color_data = 12'h332;
			{8'd108, 8'd82}: color_data = 12'hc97;
			{8'd108, 8'd83}: color_data = 12'ha86;
			{8'd108, 8'd84}: color_data = 12'h911;
			{8'd108, 8'd85}: color_data = 12'hf12;
			{8'd108, 8'd86}: color_data = 12'hf12;
			{8'd108, 8'd87}: color_data = 12'hc11;
			{8'd108, 8'd88}: color_data = 12'h944;
			{8'd108, 8'd89}: color_data = 12'h988;
			{8'd108, 8'd90}: color_data = 12'hbaa;
			{8'd108, 8'd91}: color_data = 12'hcbb;
			{8'd108, 8'd92}: color_data = 12'hccc;
			{8'd108, 8'd93}: color_data = 12'hbbb;
			{8'd108, 8'd94}: color_data = 12'hb99;
			{8'd108, 8'd95}: color_data = 12'ha77;
			{8'd108, 8'd96}: color_data = 12'h945;
			{8'd108, 8'd97}: color_data = 12'ha22;
			{8'd108, 8'd98}: color_data = 12'hd11;
			{8'd108, 8'd99}: color_data = 12'he12;
			{8'd108, 8'd100}: color_data = 12'h843;
			{8'd108, 8'd101}: color_data = 12'hc97;
			{8'd108, 8'd102}: color_data = 12'hc97;
			{8'd108, 8'd103}: color_data = 12'hb86;
			{8'd108, 8'd104}: color_data = 12'h864;
			{8'd108, 8'd105}: color_data = 12'hc97;
			{8'd108, 8'd106}: color_data = 12'hc97;
			{8'd108, 8'd107}: color_data = 12'hc97;
			{8'd108, 8'd108}: color_data = 12'hc97;
			{8'd108, 8'd109}: color_data = 12'hc97;
			{8'd108, 8'd110}: color_data = 12'hc97;
			{8'd108, 8'd111}: color_data = 12'hc97;
			{8'd108, 8'd112}: color_data = 12'hc97;
			{8'd108, 8'd113}: color_data = 12'hc97;
			{8'd108, 8'd114}: color_data = 12'hc97;
			{8'd108, 8'd115}: color_data = 12'hc97;
			{8'd108, 8'd116}: color_data = 12'hc97;
			{8'd108, 8'd117}: color_data = 12'hc97;
			{8'd108, 8'd118}: color_data = 12'hc97;
			{8'd108, 8'd119}: color_data = 12'hc97;
			{8'd108, 8'd120}: color_data = 12'hc97;
			{8'd108, 8'd121}: color_data = 12'hc97;
			{8'd108, 8'd122}: color_data = 12'hc97;
			{8'd108, 8'd123}: color_data = 12'hc97;
			{8'd108, 8'd124}: color_data = 12'hc97;
			{8'd108, 8'd125}: color_data = 12'hb86;
			{8'd108, 8'd126}: color_data = 12'h975;
			{8'd108, 8'd127}: color_data = 12'h655;
			{8'd108, 8'd128}: color_data = 12'h345;
			{8'd108, 8'd129}: color_data = 12'h036;
			{8'd108, 8'd130}: color_data = 12'h048;
			{8'd108, 8'd131}: color_data = 12'h059;
			{8'd108, 8'd132}: color_data = 12'h05a;
			{8'd108, 8'd133}: color_data = 12'h05a;
			{8'd108, 8'd134}: color_data = 12'h05a;
			{8'd108, 8'd135}: color_data = 12'h059;
			{8'd108, 8'd136}: color_data = 12'h048;
			{8'd108, 8'd137}: color_data = 12'h035;
			{8'd108, 8'd138}: color_data = 12'h001;
			{8'd108, 8'd139}: color_data = 12'h000;
			{8'd108, 8'd147}: color_data = 12'h000;
			{8'd108, 8'd148}: color_data = 12'h521;
			{8'd108, 8'd149}: color_data = 12'h843;
			{8'd108, 8'd150}: color_data = 12'h842;
			{8'd108, 8'd151}: color_data = 12'h842;
			{8'd108, 8'd152}: color_data = 12'h842;
			{8'd108, 8'd153}: color_data = 12'h842;
			{8'd108, 8'd154}: color_data = 12'h842;
			{8'd108, 8'd155}: color_data = 12'h842;
			{8'd108, 8'd156}: color_data = 12'h842;
			{8'd108, 8'd157}: color_data = 12'h753;
			{8'd108, 8'd158}: color_data = 12'h532;
			{8'd109, 8'd3}: color_data = 12'hfc5;
			{8'd109, 8'd4}: color_data = 12'hfc5;
			{8'd109, 8'd5}: color_data = 12'hfc5;
			{8'd109, 8'd6}: color_data = 12'hfc4;
			{8'd109, 8'd7}: color_data = 12'hfc5;
			{8'd109, 8'd8}: color_data = 12'hfd7;
			{8'd109, 8'd9}: color_data = 12'hea2;
			{8'd109, 8'd10}: color_data = 12'hd90;
			{8'd109, 8'd11}: color_data = 12'hd90;
			{8'd109, 8'd12}: color_data = 12'hd90;
			{8'd109, 8'd13}: color_data = 12'hd90;
			{8'd109, 8'd14}: color_data = 12'hd90;
			{8'd109, 8'd15}: color_data = 12'hd90;
			{8'd109, 8'd16}: color_data = 12'hd90;
			{8'd109, 8'd17}: color_data = 12'hfb3;
			{8'd109, 8'd18}: color_data = 12'hfc5;
			{8'd109, 8'd19}: color_data = 12'hfc5;
			{8'd109, 8'd47}: color_data = 12'h400;
			{8'd109, 8'd48}: color_data = 12'hd12;
			{8'd109, 8'd49}: color_data = 12'hf12;
			{8'd109, 8'd50}: color_data = 12'hb11;
			{8'd109, 8'd51}: color_data = 12'h200;
			{8'd109, 8'd53}: color_data = 12'h000;
			{8'd109, 8'd54}: color_data = 12'h652;
			{8'd109, 8'd55}: color_data = 12'hb94;
			{8'd109, 8'd56}: color_data = 12'hdb6;
			{8'd109, 8'd57}: color_data = 12'hb95;
			{8'd109, 8'd58}: color_data = 12'h873;
			{8'd109, 8'd59}: color_data = 12'h873;
			{8'd109, 8'd60}: color_data = 12'h873;
			{8'd109, 8'd61}: color_data = 12'h875;
			{8'd109, 8'd62}: color_data = 12'hfca;
			{8'd109, 8'd63}: color_data = 12'hfdb;
			{8'd109, 8'd64}: color_data = 12'hfda;
			{8'd109, 8'd65}: color_data = 12'hfda;
			{8'd109, 8'd66}: color_data = 12'hfda;
			{8'd109, 8'd67}: color_data = 12'hfda;
			{8'd109, 8'd68}: color_data = 12'hfda;
			{8'd109, 8'd69}: color_data = 12'hfda;
			{8'd109, 8'd70}: color_data = 12'hfdb;
			{8'd109, 8'd71}: color_data = 12'h543;
			{8'd109, 8'd72}: color_data = 12'h000;
			{8'd109, 8'd73}: color_data = 12'h000;
			{8'd109, 8'd74}: color_data = 12'h000;
			{8'd109, 8'd75}: color_data = 12'h000;
			{8'd109, 8'd76}: color_data = 12'h765;
			{8'd109, 8'd77}: color_data = 12'ha86;
			{8'd109, 8'd78}: color_data = 12'h543;
			{8'd109, 8'd79}: color_data = 12'h012;
			{8'd109, 8'd80}: color_data = 12'h333;
			{8'd109, 8'd81}: color_data = 12'h975;
			{8'd109, 8'd82}: color_data = 12'h975;
			{8'd109, 8'd83}: color_data = 12'ha76;
			{8'd109, 8'd84}: color_data = 12'h632;
			{8'd109, 8'd85}: color_data = 12'hc11;
			{8'd109, 8'd86}: color_data = 12'hf12;
			{8'd109, 8'd87}: color_data = 12'hf12;
			{8'd109, 8'd88}: color_data = 12'hd11;
			{8'd109, 8'd89}: color_data = 12'h901;
			{8'd109, 8'd90}: color_data = 12'hd11;
			{8'd109, 8'd91}: color_data = 12'hc11;
			{8'd109, 8'd92}: color_data = 12'hc11;
			{8'd109, 8'd93}: color_data = 12'hc11;
			{8'd109, 8'd94}: color_data = 12'hd11;
			{8'd109, 8'd95}: color_data = 12'he11;
			{8'd109, 8'd96}: color_data = 12'he11;
			{8'd109, 8'd97}: color_data = 12'hf12;
			{8'd109, 8'd98}: color_data = 12'hf12;
			{8'd109, 8'd99}: color_data = 12'hf12;
			{8'd109, 8'd100}: color_data = 12'h922;
			{8'd109, 8'd101}: color_data = 12'hb87;
			{8'd109, 8'd102}: color_data = 12'hc97;
			{8'd109, 8'd103}: color_data = 12'hc97;
			{8'd109, 8'd104}: color_data = 12'h865;
			{8'd109, 8'd105}: color_data = 12'ha76;
			{8'd109, 8'd106}: color_data = 12'hc97;
			{8'd109, 8'd107}: color_data = 12'hc97;
			{8'd109, 8'd108}: color_data = 12'hc97;
			{8'd109, 8'd109}: color_data = 12'hc97;
			{8'd109, 8'd110}: color_data = 12'hc97;
			{8'd109, 8'd111}: color_data = 12'hc97;
			{8'd109, 8'd112}: color_data = 12'hc97;
			{8'd109, 8'd113}: color_data = 12'hc97;
			{8'd109, 8'd114}: color_data = 12'hc97;
			{8'd109, 8'd115}: color_data = 12'hc97;
			{8'd109, 8'd116}: color_data = 12'hc97;
			{8'd109, 8'd117}: color_data = 12'hc97;
			{8'd109, 8'd118}: color_data = 12'hc97;
			{8'd109, 8'd119}: color_data = 12'hc97;
			{8'd109, 8'd120}: color_data = 12'hc97;
			{8'd109, 8'd121}: color_data = 12'hc97;
			{8'd109, 8'd122}: color_data = 12'hc97;
			{8'd109, 8'd123}: color_data = 12'hc97;
			{8'd109, 8'd124}: color_data = 12'hc97;
			{8'd109, 8'd125}: color_data = 12'hc97;
			{8'd109, 8'd126}: color_data = 12'hc97;
			{8'd109, 8'd127}: color_data = 12'hd97;
			{8'd109, 8'd128}: color_data = 12'ha75;
			{8'd109, 8'd129}: color_data = 12'h000;
			{8'd109, 8'd130}: color_data = 12'h000;
			{8'd109, 8'd131}: color_data = 12'h000;
			{8'd109, 8'd132}: color_data = 12'h012;
			{8'd109, 8'd133}: color_data = 12'h012;
			{8'd109, 8'd134}: color_data = 12'h012;
			{8'd109, 8'd135}: color_data = 12'h001;
			{8'd109, 8'd136}: color_data = 12'h000;
			{8'd109, 8'd137}: color_data = 12'h000;
			{8'd109, 8'd148}: color_data = 12'h210;
			{8'd109, 8'd149}: color_data = 12'h842;
			{8'd109, 8'd150}: color_data = 12'h843;
			{8'd109, 8'd151}: color_data = 12'h842;
			{8'd109, 8'd152}: color_data = 12'h842;
			{8'd109, 8'd153}: color_data = 12'h842;
			{8'd109, 8'd154}: color_data = 12'h842;
			{8'd109, 8'd155}: color_data = 12'h843;
			{8'd109, 8'd156}: color_data = 12'h742;
			{8'd109, 8'd157}: color_data = 12'h642;
			{8'd109, 8'd158}: color_data = 12'h000;
			{8'd110, 8'd3}: color_data = 12'hfb5;
			{8'd110, 8'd4}: color_data = 12'hfc4;
			{8'd110, 8'd5}: color_data = 12'hfc5;
			{8'd110, 8'd6}: color_data = 12'hfc5;
			{8'd110, 8'd7}: color_data = 12'hfc4;
			{8'd110, 8'd8}: color_data = 12'hfc5;
			{8'd110, 8'd9}: color_data = 12'hea1;
			{8'd110, 8'd10}: color_data = 12'hd90;
			{8'd110, 8'd11}: color_data = 12'hd90;
			{8'd110, 8'd12}: color_data = 12'hd90;
			{8'd110, 8'd13}: color_data = 12'hd90;
			{8'd110, 8'd14}: color_data = 12'hd90;
			{8'd110, 8'd15}: color_data = 12'hd90;
			{8'd110, 8'd16}: color_data = 12'hea0;
			{8'd110, 8'd17}: color_data = 12'hfc5;
			{8'd110, 8'd18}: color_data = 12'hfc5;
			{8'd110, 8'd19}: color_data = 12'hfc6;
			{8'd110, 8'd46}: color_data = 12'h000;
			{8'd110, 8'd47}: color_data = 12'h911;
			{8'd110, 8'd48}: color_data = 12'hf12;
			{8'd110, 8'd49}: color_data = 12'hd12;
			{8'd110, 8'd50}: color_data = 12'h400;
			{8'd110, 8'd53}: color_data = 12'h000;
			{8'd110, 8'd54}: color_data = 12'h763;
			{8'd110, 8'd55}: color_data = 12'ha94;
			{8'd110, 8'd56}: color_data = 12'h763;
			{8'd110, 8'd57}: color_data = 12'hca5;
			{8'd110, 8'd58}: color_data = 12'hec6;
			{8'd110, 8'd59}: color_data = 12'hec6;
			{8'd110, 8'd60}: color_data = 12'h875;
			{8'd110, 8'd61}: color_data = 12'hfca;
			{8'd110, 8'd62}: color_data = 12'hfdb;
			{8'd110, 8'd63}: color_data = 12'hfda;
			{8'd110, 8'd64}: color_data = 12'hfda;
			{8'd110, 8'd65}: color_data = 12'hfda;
			{8'd110, 8'd66}: color_data = 12'hfda;
			{8'd110, 8'd67}: color_data = 12'hfda;
			{8'd110, 8'd68}: color_data = 12'hfda;
			{8'd110, 8'd69}: color_data = 12'hfda;
			{8'd110, 8'd70}: color_data = 12'hfdb;
			{8'd110, 8'd71}: color_data = 12'hb97;
			{8'd110, 8'd72}: color_data = 12'h000;
			{8'd110, 8'd73}: color_data = 12'h000;
			{8'd110, 8'd74}: color_data = 12'h000;
			{8'd110, 8'd75}: color_data = 12'h000;
			{8'd110, 8'd76}: color_data = 12'h965;
			{8'd110, 8'd77}: color_data = 12'hc97;
			{8'd110, 8'd78}: color_data = 12'h222;
			{8'd110, 8'd79}: color_data = 12'h112;
			{8'd110, 8'd80}: color_data = 12'h865;
			{8'd110, 8'd81}: color_data = 12'hd97;
			{8'd110, 8'd82}: color_data = 12'h864;
			{8'd110, 8'd83}: color_data = 12'h865;
			{8'd110, 8'd84}: color_data = 12'ha86;
			{8'd110, 8'd85}: color_data = 12'h844;
			{8'd110, 8'd86}: color_data = 12'hc11;
			{8'd110, 8'd87}: color_data = 12'hf12;
			{8'd110, 8'd88}: color_data = 12'hc11;
			{8'd110, 8'd89}: color_data = 12'hb11;
			{8'd110, 8'd90}: color_data = 12'hf12;
			{8'd110, 8'd91}: color_data = 12'hf12;
			{8'd110, 8'd92}: color_data = 12'hf12;
			{8'd110, 8'd93}: color_data = 12'hf12;
			{8'd110, 8'd94}: color_data = 12'hf12;
			{8'd110, 8'd95}: color_data = 12'he12;
			{8'd110, 8'd96}: color_data = 12'he12;
			{8'd110, 8'd97}: color_data = 12'he12;
			{8'd110, 8'd98}: color_data = 12'he12;
			{8'd110, 8'd99}: color_data = 12'hf12;
			{8'd110, 8'd100}: color_data = 12'hc11;
			{8'd110, 8'd101}: color_data = 12'h965;
			{8'd110, 8'd102}: color_data = 12'hc97;
			{8'd110, 8'd103}: color_data = 12'hc97;
			{8'd110, 8'd104}: color_data = 12'hc97;
			{8'd110, 8'd105}: color_data = 12'h754;
			{8'd110, 8'd106}: color_data = 12'hc97;
			{8'd110, 8'd107}: color_data = 12'hc97;
			{8'd110, 8'd108}: color_data = 12'hc97;
			{8'd110, 8'd109}: color_data = 12'hc97;
			{8'd110, 8'd110}: color_data = 12'hc97;
			{8'd110, 8'd111}: color_data = 12'hc97;
			{8'd110, 8'd112}: color_data = 12'hc97;
			{8'd110, 8'd113}: color_data = 12'hc97;
			{8'd110, 8'd114}: color_data = 12'hc97;
			{8'd110, 8'd115}: color_data = 12'hc97;
			{8'd110, 8'd116}: color_data = 12'hc97;
			{8'd110, 8'd117}: color_data = 12'hc97;
			{8'd110, 8'd118}: color_data = 12'hc97;
			{8'd110, 8'd119}: color_data = 12'hc97;
			{8'd110, 8'd120}: color_data = 12'hc97;
			{8'd110, 8'd121}: color_data = 12'hc97;
			{8'd110, 8'd122}: color_data = 12'hc97;
			{8'd110, 8'd123}: color_data = 12'hc97;
			{8'd110, 8'd124}: color_data = 12'hc97;
			{8'd110, 8'd125}: color_data = 12'hc97;
			{8'd110, 8'd126}: color_data = 12'hc97;
			{8'd110, 8'd127}: color_data = 12'hc97;
			{8'd110, 8'd128}: color_data = 12'h976;
			{8'd110, 8'd129}: color_data = 12'h000;
			{8'd110, 8'd148}: color_data = 12'h000;
			{8'd110, 8'd149}: color_data = 12'h521;
			{8'd110, 8'd150}: color_data = 12'h853;
			{8'd110, 8'd151}: color_data = 12'h842;
			{8'd110, 8'd152}: color_data = 12'h842;
			{8'd110, 8'd153}: color_data = 12'h842;
			{8'd110, 8'd154}: color_data = 12'h843;
			{8'd110, 8'd155}: color_data = 12'h742;
			{8'd110, 8'd156}: color_data = 12'h532;
			{8'd110, 8'd157}: color_data = 12'h321;
			{8'd111, 8'd2}: color_data = 12'hfd5;
			{8'd111, 8'd3}: color_data = 12'hfc5;
			{8'd111, 8'd4}: color_data = 12'hfc5;
			{8'd111, 8'd5}: color_data = 12'hfb4;
			{8'd111, 8'd6}: color_data = 12'hea0;
			{8'd111, 8'd7}: color_data = 12'hd90;
			{8'd111, 8'd8}: color_data = 12'hd90;
			{8'd111, 8'd9}: color_data = 12'hd90;
			{8'd111, 8'd10}: color_data = 12'hd90;
			{8'd111, 8'd11}: color_data = 12'hd90;
			{8'd111, 8'd12}: color_data = 12'hd90;
			{8'd111, 8'd13}: color_data = 12'heb2;
			{8'd111, 8'd14}: color_data = 12'hea2;
			{8'd111, 8'd15}: color_data = 12'hea0;
			{8'd111, 8'd16}: color_data = 12'heb2;
			{8'd111, 8'd17}: color_data = 12'hfc5;
			{8'd111, 8'd18}: color_data = 12'hfc5;
			{8'd111, 8'd46}: color_data = 12'h400;
			{8'd111, 8'd47}: color_data = 12'he12;
			{8'd111, 8'd48}: color_data = 12'hd12;
			{8'd111, 8'd49}: color_data = 12'h400;
			{8'd111, 8'd50}: color_data = 12'h000;
			{8'd111, 8'd53}: color_data = 12'h000;
			{8'd111, 8'd54}: color_data = 12'h652;
			{8'd111, 8'd55}: color_data = 12'ha94;
			{8'd111, 8'd56}: color_data = 12'hfd6;
			{8'd111, 8'd57}: color_data = 12'hfd7;
			{8'd111, 8'd58}: color_data = 12'hfe7;
			{8'd111, 8'd59}: color_data = 12'hca5;
			{8'd111, 8'd60}: color_data = 12'hca8;
			{8'd111, 8'd61}: color_data = 12'hfdb;
			{8'd111, 8'd62}: color_data = 12'hfda;
			{8'd111, 8'd63}: color_data = 12'hfda;
			{8'd111, 8'd64}: color_data = 12'hfda;
			{8'd111, 8'd65}: color_data = 12'hfda;
			{8'd111, 8'd66}: color_data = 12'hfda;
			{8'd111, 8'd67}: color_data = 12'hfda;
			{8'd111, 8'd68}: color_data = 12'hfda;
			{8'd111, 8'd69}: color_data = 12'hfda;
			{8'd111, 8'd70}: color_data = 12'hfdb;
			{8'd111, 8'd71}: color_data = 12'heb9;
			{8'd111, 8'd72}: color_data = 12'h100;
			{8'd111, 8'd73}: color_data = 12'h000;
			{8'd111, 8'd74}: color_data = 12'h111;
			{8'd111, 8'd75}: color_data = 12'h975;
			{8'd111, 8'd76}: color_data = 12'hda8;
			{8'd111, 8'd77}: color_data = 12'h975;
			{8'd111, 8'd78}: color_data = 12'h012;
			{8'd111, 8'd79}: color_data = 12'h223;
			{8'd111, 8'd80}: color_data = 12'hc97;
			{8'd111, 8'd81}: color_data = 12'hc97;
			{8'd111, 8'd82}: color_data = 12'hb87;
			{8'd111, 8'd83}: color_data = 12'h643;
			{8'd111, 8'd84}: color_data = 12'hb86;
			{8'd111, 8'd85}: color_data = 12'hc97;
			{8'd111, 8'd86}: color_data = 12'h843;
			{8'd111, 8'd87}: color_data = 12'hd11;
			{8'd111, 8'd88}: color_data = 12'hc11;
			{8'd111, 8'd89}: color_data = 12'hb11;
			{8'd111, 8'd90}: color_data = 12'hf12;
			{8'd111, 8'd91}: color_data = 12'he12;
			{8'd111, 8'd92}: color_data = 12'he12;
			{8'd111, 8'd93}: color_data = 12'he12;
			{8'd111, 8'd94}: color_data = 12'he12;
			{8'd111, 8'd95}: color_data = 12'he12;
			{8'd111, 8'd96}: color_data = 12'he12;
			{8'd111, 8'd97}: color_data = 12'he12;
			{8'd111, 8'd98}: color_data = 12'he12;
			{8'd111, 8'd99}: color_data = 12'he12;
			{8'd111, 8'd100}: color_data = 12'he12;
			{8'd111, 8'd101}: color_data = 12'h843;
			{8'd111, 8'd102}: color_data = 12'hc97;
			{8'd111, 8'd103}: color_data = 12'hc97;
			{8'd111, 8'd104}: color_data = 12'hc97;
			{8'd111, 8'd105}: color_data = 12'ha86;
			{8'd111, 8'd106}: color_data = 12'ha86;
			{8'd111, 8'd107}: color_data = 12'hc97;
			{8'd111, 8'd108}: color_data = 12'hc97;
			{8'd111, 8'd109}: color_data = 12'hc97;
			{8'd111, 8'd110}: color_data = 12'hc97;
			{8'd111, 8'd111}: color_data = 12'hc97;
			{8'd111, 8'd112}: color_data = 12'hc97;
			{8'd111, 8'd113}: color_data = 12'hc97;
			{8'd111, 8'd114}: color_data = 12'hc97;
			{8'd111, 8'd115}: color_data = 12'hc97;
			{8'd111, 8'd116}: color_data = 12'hc97;
			{8'd111, 8'd117}: color_data = 12'hc97;
			{8'd111, 8'd118}: color_data = 12'hc97;
			{8'd111, 8'd119}: color_data = 12'hc97;
			{8'd111, 8'd120}: color_data = 12'hc97;
			{8'd111, 8'd121}: color_data = 12'hc97;
			{8'd111, 8'd122}: color_data = 12'hc97;
			{8'd111, 8'd123}: color_data = 12'hc97;
			{8'd111, 8'd124}: color_data = 12'hc97;
			{8'd111, 8'd125}: color_data = 12'hc97;
			{8'd111, 8'd126}: color_data = 12'hc97;
			{8'd111, 8'd127}: color_data = 12'hc97;
			{8'd111, 8'd128}: color_data = 12'h975;
			{8'd111, 8'd129}: color_data = 12'h000;
			{8'd111, 8'd149}: color_data = 12'h100;
			{8'd111, 8'd150}: color_data = 12'h732;
			{8'd111, 8'd151}: color_data = 12'h843;
			{8'd111, 8'd152}: color_data = 12'h842;
			{8'd111, 8'd153}: color_data = 12'h843;
			{8'd111, 8'd154}: color_data = 12'h842;
			{8'd111, 8'd155}: color_data = 12'h321;
			{8'd111, 8'd156}: color_data = 12'h210;
			{8'd112, 8'd1}: color_data = 12'heb5;
			{8'd112, 8'd2}: color_data = 12'hfc5;
			{8'd112, 8'd3}: color_data = 12'hfc5;
			{8'd112, 8'd4}: color_data = 12'hfc4;
			{8'd112, 8'd5}: color_data = 12'hda0;
			{8'd112, 8'd6}: color_data = 12'hd90;
			{8'd112, 8'd7}: color_data = 12'hd90;
			{8'd112, 8'd8}: color_data = 12'hd90;
			{8'd112, 8'd9}: color_data = 12'hd90;
			{8'd112, 8'd10}: color_data = 12'hd90;
			{8'd112, 8'd11}: color_data = 12'hd90;
			{8'd112, 8'd12}: color_data = 12'hd90;
			{8'd112, 8'd13}: color_data = 12'hfb4;
			{8'd112, 8'd14}: color_data = 12'hfd7;
			{8'd112, 8'd15}: color_data = 12'hfc5;
			{8'd112, 8'd16}: color_data = 12'hfc5;
			{8'd112, 8'd17}: color_data = 12'hfc5;
			{8'd112, 8'd18}: color_data = 12'hfc5;
			{8'd112, 8'd45}: color_data = 12'h000;
			{8'd112, 8'd46}: color_data = 12'ha11;
			{8'd112, 8'd47}: color_data = 12'hc11;
			{8'd112, 8'd48}: color_data = 12'h400;
			{8'd112, 8'd49}: color_data = 12'h000;
			{8'd112, 8'd54}: color_data = 12'h431;
			{8'd112, 8'd55}: color_data = 12'hec6;
			{8'd112, 8'd56}: color_data = 12'hfd7;
			{8'd112, 8'd57}: color_data = 12'hfe7;
			{8'd112, 8'd58}: color_data = 12'hfe7;
			{8'd112, 8'd59}: color_data = 12'ha84;
			{8'd112, 8'd60}: color_data = 12'hdb9;
			{8'd112, 8'd61}: color_data = 12'hfdb;
			{8'd112, 8'd62}: color_data = 12'hfda;
			{8'd112, 8'd63}: color_data = 12'hfda;
			{8'd112, 8'd64}: color_data = 12'hfda;
			{8'd112, 8'd65}: color_data = 12'hfda;
			{8'd112, 8'd66}: color_data = 12'hfda;
			{8'd112, 8'd67}: color_data = 12'hfda;
			{8'd112, 8'd68}: color_data = 12'hfda;
			{8'd112, 8'd69}: color_data = 12'hfda;
			{8'd112, 8'd70}: color_data = 12'hfdb;
			{8'd112, 8'd71}: color_data = 12'heca;
			{8'd112, 8'd72}: color_data = 12'h110;
			{8'd112, 8'd73}: color_data = 12'h000;
			{8'd112, 8'd74}: color_data = 12'h432;
			{8'd112, 8'd75}: color_data = 12'hda8;
			{8'd112, 8'd76}: color_data = 12'hc97;
			{8'd112, 8'd77}: color_data = 12'h644;
			{8'd112, 8'd78}: color_data = 12'h012;
			{8'd112, 8'd79}: color_data = 12'h544;
			{8'd112, 8'd80}: color_data = 12'hc97;
			{8'd112, 8'd81}: color_data = 12'hc97;
			{8'd112, 8'd82}: color_data = 12'hc97;
			{8'd112, 8'd83}: color_data = 12'hb87;
			{8'd112, 8'd84}: color_data = 12'h754;
			{8'd112, 8'd85}: color_data = 12'h865;
			{8'd112, 8'd86}: color_data = 12'h865;
			{8'd112, 8'd87}: color_data = 12'h622;
			{8'd112, 8'd88}: color_data = 12'hb11;
			{8'd112, 8'd89}: color_data = 12'hb11;
			{8'd112, 8'd90}: color_data = 12'hf12;
			{8'd112, 8'd91}: color_data = 12'he12;
			{8'd112, 8'd92}: color_data = 12'he12;
			{8'd112, 8'd93}: color_data = 12'he12;
			{8'd112, 8'd94}: color_data = 12'he12;
			{8'd112, 8'd95}: color_data = 12'he12;
			{8'd112, 8'd96}: color_data = 12'he12;
			{8'd112, 8'd97}: color_data = 12'he12;
			{8'd112, 8'd98}: color_data = 12'he12;
			{8'd112, 8'd99}: color_data = 12'he12;
			{8'd112, 8'd100}: color_data = 12'hf12;
			{8'd112, 8'd101}: color_data = 12'h832;
			{8'd112, 8'd102}: color_data = 12'hc97;
			{8'd112, 8'd103}: color_data = 12'hc97;
			{8'd112, 8'd104}: color_data = 12'hc97;
			{8'd112, 8'd105}: color_data = 12'hc97;
			{8'd112, 8'd106}: color_data = 12'hc97;
			{8'd112, 8'd107}: color_data = 12'hc97;
			{8'd112, 8'd108}: color_data = 12'hc97;
			{8'd112, 8'd109}: color_data = 12'hc97;
			{8'd112, 8'd110}: color_data = 12'hc97;
			{8'd112, 8'd111}: color_data = 12'hc97;
			{8'd112, 8'd112}: color_data = 12'hc97;
			{8'd112, 8'd113}: color_data = 12'hc97;
			{8'd112, 8'd114}: color_data = 12'hc97;
			{8'd112, 8'd115}: color_data = 12'hc97;
			{8'd112, 8'd116}: color_data = 12'hc97;
			{8'd112, 8'd117}: color_data = 12'hc97;
			{8'd112, 8'd118}: color_data = 12'hc97;
			{8'd112, 8'd119}: color_data = 12'hc97;
			{8'd112, 8'd120}: color_data = 12'hc97;
			{8'd112, 8'd121}: color_data = 12'hc97;
			{8'd112, 8'd122}: color_data = 12'hc97;
			{8'd112, 8'd123}: color_data = 12'hc97;
			{8'd112, 8'd124}: color_data = 12'hc97;
			{8'd112, 8'd125}: color_data = 12'hc97;
			{8'd112, 8'd126}: color_data = 12'hc97;
			{8'd112, 8'd127}: color_data = 12'hc97;
			{8'd112, 8'd128}: color_data = 12'h975;
			{8'd112, 8'd129}: color_data = 12'h000;
			{8'd112, 8'd150}: color_data = 12'h210;
			{8'd112, 8'd151}: color_data = 12'h632;
			{8'd112, 8'd152}: color_data = 12'h842;
			{8'd112, 8'd153}: color_data = 12'h842;
			{8'd112, 8'd154}: color_data = 12'h421;
			{8'd112, 8'd155}: color_data = 12'h000;
			{8'd113, 8'd1}: color_data = 12'hfc5;
			{8'd113, 8'd2}: color_data = 12'hfc5;
			{8'd113, 8'd3}: color_data = 12'hfc4;
			{8'd113, 8'd4}: color_data = 12'hea0;
			{8'd113, 8'd5}: color_data = 12'hd90;
			{8'd113, 8'd6}: color_data = 12'hd90;
			{8'd113, 8'd7}: color_data = 12'hd90;
			{8'd113, 8'd8}: color_data = 12'hd90;
			{8'd113, 8'd9}: color_data = 12'hd90;
			{8'd113, 8'd10}: color_data = 12'hd90;
			{8'd113, 8'd11}: color_data = 12'hd90;
			{8'd113, 8'd12}: color_data = 12'hd90;
			{8'd113, 8'd13}: color_data = 12'hea0;
			{8'd113, 8'd14}: color_data = 12'hfc5;
			{8'd113, 8'd15}: color_data = 12'hfc5;
			{8'd113, 8'd16}: color_data = 12'hfc5;
			{8'd113, 8'd17}: color_data = 12'hfc5;
			{8'd113, 8'd18}: color_data = 12'hf0f;
			{8'd113, 8'd45}: color_data = 12'h400;
			{8'd113, 8'd46}: color_data = 12'h811;
			{8'd113, 8'd47}: color_data = 12'h200;
			{8'd113, 8'd54}: color_data = 12'h000;
			{8'd113, 8'd55}: color_data = 12'h221;
			{8'd113, 8'd56}: color_data = 12'h652;
			{8'd113, 8'd57}: color_data = 12'h973;
			{8'd113, 8'd58}: color_data = 12'h873;
			{8'd113, 8'd59}: color_data = 12'h652;
			{8'd113, 8'd60}: color_data = 12'hdb9;
			{8'd113, 8'd61}: color_data = 12'hfdb;
			{8'd113, 8'd62}: color_data = 12'hfda;
			{8'd113, 8'd63}: color_data = 12'hfda;
			{8'd113, 8'd64}: color_data = 12'hfda;
			{8'd113, 8'd65}: color_data = 12'hfda;
			{8'd113, 8'd66}: color_data = 12'hfda;
			{8'd113, 8'd67}: color_data = 12'hfda;
			{8'd113, 8'd68}: color_data = 12'hfda;
			{8'd113, 8'd69}: color_data = 12'hfda;
			{8'd113, 8'd70}: color_data = 12'hfdb;
			{8'd113, 8'd71}: color_data = 12'hca8;
			{8'd113, 8'd72}: color_data = 12'h000;
			{8'd113, 8'd73}: color_data = 12'h000;
			{8'd113, 8'd74}: color_data = 12'h543;
			{8'd113, 8'd75}: color_data = 12'hd97;
			{8'd113, 8'd76}: color_data = 12'hc97;
			{8'd113, 8'd77}: color_data = 12'h323;
			{8'd113, 8'd78}: color_data = 12'h012;
			{8'd113, 8'd79}: color_data = 12'h865;
			{8'd113, 8'd80}: color_data = 12'hc97;
			{8'd113, 8'd81}: color_data = 12'hc97;
			{8'd113, 8'd82}: color_data = 12'hc97;
			{8'd113, 8'd83}: color_data = 12'hc97;
			{8'd113, 8'd84}: color_data = 12'hc97;
			{8'd113, 8'd85}: color_data = 12'hb86;
			{8'd113, 8'd86}: color_data = 12'hb86;
			{8'd113, 8'd87}: color_data = 12'hb86;
			{8'd113, 8'd88}: color_data = 12'h622;
			{8'd113, 8'd89}: color_data = 12'ha11;
			{8'd113, 8'd90}: color_data = 12'hf12;
			{8'd113, 8'd91}: color_data = 12'he12;
			{8'd113, 8'd92}: color_data = 12'he12;
			{8'd113, 8'd93}: color_data = 12'he12;
			{8'd113, 8'd94}: color_data = 12'he12;
			{8'd113, 8'd95}: color_data = 12'he12;
			{8'd113, 8'd96}: color_data = 12'he12;
			{8'd113, 8'd97}: color_data = 12'he12;
			{8'd113, 8'd98}: color_data = 12'he12;
			{8'd113, 8'd99}: color_data = 12'he12;
			{8'd113, 8'd100}: color_data = 12'hf12;
			{8'd113, 8'd101}: color_data = 12'h922;
			{8'd113, 8'd102}: color_data = 12'hb97;
			{8'd113, 8'd103}: color_data = 12'hc97;
			{8'd113, 8'd104}: color_data = 12'hc97;
			{8'd113, 8'd105}: color_data = 12'hc97;
			{8'd113, 8'd106}: color_data = 12'hc97;
			{8'd113, 8'd107}: color_data = 12'hc97;
			{8'd113, 8'd108}: color_data = 12'hc97;
			{8'd113, 8'd109}: color_data = 12'hc97;
			{8'd113, 8'd110}: color_data = 12'hc97;
			{8'd113, 8'd111}: color_data = 12'hc97;
			{8'd113, 8'd112}: color_data = 12'hc97;
			{8'd113, 8'd113}: color_data = 12'hc97;
			{8'd113, 8'd114}: color_data = 12'hc97;
			{8'd113, 8'd115}: color_data = 12'hc97;
			{8'd113, 8'd116}: color_data = 12'hc97;
			{8'd113, 8'd117}: color_data = 12'hc97;
			{8'd113, 8'd118}: color_data = 12'hc97;
			{8'd113, 8'd119}: color_data = 12'hc97;
			{8'd113, 8'd120}: color_data = 12'hc97;
			{8'd113, 8'd121}: color_data = 12'hc97;
			{8'd113, 8'd122}: color_data = 12'hc97;
			{8'd113, 8'd123}: color_data = 12'hc97;
			{8'd113, 8'd124}: color_data = 12'hc97;
			{8'd113, 8'd125}: color_data = 12'hc97;
			{8'd113, 8'd126}: color_data = 12'hc97;
			{8'd113, 8'd127}: color_data = 12'hc97;
			{8'd113, 8'd128}: color_data = 12'h965;
			{8'd113, 8'd129}: color_data = 12'h000;
			{8'd113, 8'd150}: color_data = 12'h000;
			{8'd113, 8'd151}: color_data = 12'h000;
			{8'd113, 8'd152}: color_data = 12'h210;
			{8'd113, 8'd153}: color_data = 12'h210;
			{8'd113, 8'd154}: color_data = 12'h000;
			{8'd114, 8'd0}: color_data = 12'hfc6;
			{8'd114, 8'd1}: color_data = 12'hfc5;
			{8'd114, 8'd2}: color_data = 12'hfc5;
			{8'd114, 8'd3}: color_data = 12'hea1;
			{8'd114, 8'd4}: color_data = 12'hd90;
			{8'd114, 8'd5}: color_data = 12'hd90;
			{8'd114, 8'd6}: color_data = 12'hd90;
			{8'd114, 8'd7}: color_data = 12'hd90;
			{8'd114, 8'd8}: color_data = 12'hd90;
			{8'd114, 8'd9}: color_data = 12'hd90;
			{8'd114, 8'd10}: color_data = 12'hd90;
			{8'd114, 8'd11}: color_data = 12'hd90;
			{8'd114, 8'd12}: color_data = 12'hd90;
			{8'd114, 8'd13}: color_data = 12'hd90;
			{8'd114, 8'd14}: color_data = 12'heb2;
			{8'd114, 8'd15}: color_data = 12'hfc5;
			{8'd114, 8'd16}: color_data = 12'hfc5;
			{8'd114, 8'd17}: color_data = 12'hfd6;
			{8'd114, 8'd44}: color_data = 12'h000;
			{8'd114, 8'd45}: color_data = 12'h100;
			{8'd114, 8'd46}: color_data = 12'h200;
			{8'd114, 8'd57}: color_data = 12'h221;
			{8'd114, 8'd58}: color_data = 12'h763;
			{8'd114, 8'd59}: color_data = 12'h652;
			{8'd114, 8'd60}: color_data = 12'ha97;
			{8'd114, 8'd61}: color_data = 12'hfdb;
			{8'd114, 8'd62}: color_data = 12'hfda;
			{8'd114, 8'd63}: color_data = 12'hfda;
			{8'd114, 8'd64}: color_data = 12'hfda;
			{8'd114, 8'd65}: color_data = 12'hfda;
			{8'd114, 8'd66}: color_data = 12'hfda;
			{8'd114, 8'd67}: color_data = 12'hfda;
			{8'd114, 8'd68}: color_data = 12'hfda;
			{8'd114, 8'd69}: color_data = 12'hfda;
			{8'd114, 8'd70}: color_data = 12'hfdb;
			{8'd114, 8'd71}: color_data = 12'h654;
			{8'd114, 8'd72}: color_data = 12'h000;
			{8'd114, 8'd73}: color_data = 12'h000;
			{8'd114, 8'd74}: color_data = 12'h865;
			{8'd114, 8'd75}: color_data = 12'hd97;
			{8'd114, 8'd76}: color_data = 12'ha76;
			{8'd114, 8'd77}: color_data = 12'h112;
			{8'd114, 8'd78}: color_data = 12'h122;
			{8'd114, 8'd79}: color_data = 12'ha86;
			{8'd114, 8'd80}: color_data = 12'hc97;
			{8'd114, 8'd81}: color_data = 12'hc97;
			{8'd114, 8'd82}: color_data = 12'hc97;
			{8'd114, 8'd83}: color_data = 12'hc97;
			{8'd114, 8'd84}: color_data = 12'hc97;
			{8'd114, 8'd85}: color_data = 12'hc97;
			{8'd114, 8'd86}: color_data = 12'hc97;
			{8'd114, 8'd87}: color_data = 12'hc97;
			{8'd114, 8'd88}: color_data = 12'h975;
			{8'd114, 8'd89}: color_data = 12'h711;
			{8'd114, 8'd90}: color_data = 12'hf12;
			{8'd114, 8'd91}: color_data = 12'he12;
			{8'd114, 8'd92}: color_data = 12'he12;
			{8'd114, 8'd93}: color_data = 12'he12;
			{8'd114, 8'd94}: color_data = 12'he12;
			{8'd114, 8'd95}: color_data = 12'he12;
			{8'd114, 8'd96}: color_data = 12'he12;
			{8'd114, 8'd97}: color_data = 12'he12;
			{8'd114, 8'd98}: color_data = 12'he12;
			{8'd114, 8'd99}: color_data = 12'he12;
			{8'd114, 8'd100}: color_data = 12'hf12;
			{8'd114, 8'd101}: color_data = 12'h922;
			{8'd114, 8'd102}: color_data = 12'hb97;
			{8'd114, 8'd103}: color_data = 12'hc97;
			{8'd114, 8'd104}: color_data = 12'hc97;
			{8'd114, 8'd105}: color_data = 12'hc97;
			{8'd114, 8'd106}: color_data = 12'hc97;
			{8'd114, 8'd107}: color_data = 12'hc97;
			{8'd114, 8'd108}: color_data = 12'hc97;
			{8'd114, 8'd109}: color_data = 12'hc97;
			{8'd114, 8'd110}: color_data = 12'hc97;
			{8'd114, 8'd111}: color_data = 12'hc97;
			{8'd114, 8'd112}: color_data = 12'hc97;
			{8'd114, 8'd113}: color_data = 12'hc97;
			{8'd114, 8'd114}: color_data = 12'hc97;
			{8'd114, 8'd115}: color_data = 12'hc97;
			{8'd114, 8'd116}: color_data = 12'hc97;
			{8'd114, 8'd117}: color_data = 12'hc97;
			{8'd114, 8'd118}: color_data = 12'hc97;
			{8'd114, 8'd119}: color_data = 12'hc97;
			{8'd114, 8'd120}: color_data = 12'hc97;
			{8'd114, 8'd121}: color_data = 12'hc97;
			{8'd114, 8'd122}: color_data = 12'hc97;
			{8'd114, 8'd123}: color_data = 12'hc97;
			{8'd114, 8'd124}: color_data = 12'hc97;
			{8'd114, 8'd125}: color_data = 12'hc97;
			{8'd114, 8'd126}: color_data = 12'hc97;
			{8'd114, 8'd127}: color_data = 12'hc97;
			{8'd114, 8'd128}: color_data = 12'h865;
			{8'd114, 8'd129}: color_data = 12'h000;
			{8'd115, 8'd0}: color_data = 12'hfc5;
			{8'd115, 8'd1}: color_data = 12'hfc5;
			{8'd115, 8'd2}: color_data = 12'hfc4;
			{8'd115, 8'd3}: color_data = 12'hd90;
			{8'd115, 8'd4}: color_data = 12'hd90;
			{8'd115, 8'd5}: color_data = 12'hd90;
			{8'd115, 8'd6}: color_data = 12'hd90;
			{8'd115, 8'd7}: color_data = 12'hd90;
			{8'd115, 8'd8}: color_data = 12'hd90;
			{8'd115, 8'd9}: color_data = 12'hd90;
			{8'd115, 8'd10}: color_data = 12'hd90;
			{8'd115, 8'd11}: color_data = 12'hd90;
			{8'd115, 8'd12}: color_data = 12'hd90;
			{8'd115, 8'd13}: color_data = 12'hd90;
			{8'd115, 8'd14}: color_data = 12'hda0;
			{8'd115, 8'd15}: color_data = 12'hfc5;
			{8'd115, 8'd16}: color_data = 12'hfc5;
			{8'd115, 8'd17}: color_data = 12'hfc5;
			{8'd115, 8'd44}: color_data = 12'h000;
			{8'd115, 8'd45}: color_data = 12'h000;
			{8'd115, 8'd56}: color_data = 12'h321;
			{8'd115, 8'd57}: color_data = 12'h873;
			{8'd115, 8'd58}: color_data = 12'h984;
			{8'd115, 8'd59}: color_data = 12'h973;
			{8'd115, 8'd60}: color_data = 12'h985;
			{8'd115, 8'd61}: color_data = 12'hfdb;
			{8'd115, 8'd62}: color_data = 12'hfda;
			{8'd115, 8'd63}: color_data = 12'hfda;
			{8'd115, 8'd64}: color_data = 12'hfda;
			{8'd115, 8'd65}: color_data = 12'hfda;
			{8'd115, 8'd66}: color_data = 12'hfda;
			{8'd115, 8'd67}: color_data = 12'hfda;
			{8'd115, 8'd68}: color_data = 12'hfda;
			{8'd115, 8'd69}: color_data = 12'hfdb;
			{8'd115, 8'd70}: color_data = 12'hca8;
			{8'd115, 8'd71}: color_data = 12'h864;
			{8'd115, 8'd72}: color_data = 12'h865;
			{8'd115, 8'd73}: color_data = 12'h975;
			{8'd115, 8'd74}: color_data = 12'hc97;
			{8'd115, 8'd75}: color_data = 12'hd97;
			{8'd115, 8'd76}: color_data = 12'h754;
			{8'd115, 8'd77}: color_data = 12'h012;
			{8'd115, 8'd78}: color_data = 12'h223;
			{8'd115, 8'd79}: color_data = 12'hc97;
			{8'd115, 8'd80}: color_data = 12'hc97;
			{8'd115, 8'd81}: color_data = 12'hc97;
			{8'd115, 8'd82}: color_data = 12'hc97;
			{8'd115, 8'd83}: color_data = 12'hc97;
			{8'd115, 8'd84}: color_data = 12'hc97;
			{8'd115, 8'd85}: color_data = 12'hc97;
			{8'd115, 8'd86}: color_data = 12'hc97;
			{8'd115, 8'd87}: color_data = 12'hc97;
			{8'd115, 8'd88}: color_data = 12'hc97;
			{8'd115, 8'd89}: color_data = 12'h743;
			{8'd115, 8'd90}: color_data = 12'hd11;
			{8'd115, 8'd91}: color_data = 12'hf12;
			{8'd115, 8'd92}: color_data = 12'he12;
			{8'd115, 8'd93}: color_data = 12'he12;
			{8'd115, 8'd94}: color_data = 12'he12;
			{8'd115, 8'd95}: color_data = 12'he12;
			{8'd115, 8'd96}: color_data = 12'he12;
			{8'd115, 8'd97}: color_data = 12'he12;
			{8'd115, 8'd98}: color_data = 12'he12;
			{8'd115, 8'd99}: color_data = 12'he12;
			{8'd115, 8'd100}: color_data = 12'he12;
			{8'd115, 8'd101}: color_data = 12'h833;
			{8'd115, 8'd102}: color_data = 12'hc97;
			{8'd115, 8'd103}: color_data = 12'hc97;
			{8'd115, 8'd104}: color_data = 12'hc97;
			{8'd115, 8'd105}: color_data = 12'hc97;
			{8'd115, 8'd106}: color_data = 12'hc97;
			{8'd115, 8'd107}: color_data = 12'hc97;
			{8'd115, 8'd108}: color_data = 12'hc97;
			{8'd115, 8'd109}: color_data = 12'hc97;
			{8'd115, 8'd110}: color_data = 12'hc97;
			{8'd115, 8'd111}: color_data = 12'hc97;
			{8'd115, 8'd112}: color_data = 12'hc97;
			{8'd115, 8'd113}: color_data = 12'hc97;
			{8'd115, 8'd114}: color_data = 12'hc97;
			{8'd115, 8'd115}: color_data = 12'hc97;
			{8'd115, 8'd116}: color_data = 12'hc97;
			{8'd115, 8'd117}: color_data = 12'hc97;
			{8'd115, 8'd118}: color_data = 12'hc97;
			{8'd115, 8'd119}: color_data = 12'hc97;
			{8'd115, 8'd120}: color_data = 12'hc97;
			{8'd115, 8'd121}: color_data = 12'hc97;
			{8'd115, 8'd122}: color_data = 12'hc97;
			{8'd115, 8'd123}: color_data = 12'hc97;
			{8'd115, 8'd124}: color_data = 12'hc97;
			{8'd115, 8'd125}: color_data = 12'hc97;
			{8'd115, 8'd126}: color_data = 12'hc97;
			{8'd115, 8'd127}: color_data = 12'hd97;
			{8'd115, 8'd128}: color_data = 12'h865;
			{8'd115, 8'd129}: color_data = 12'h000;
			{8'd116, 8'd0}: color_data = 12'hfc4;
			{8'd116, 8'd1}: color_data = 12'hfc5;
			{8'd116, 8'd2}: color_data = 12'hfb3;
			{8'd116, 8'd3}: color_data = 12'hd90;
			{8'd116, 8'd4}: color_data = 12'hd90;
			{8'd116, 8'd5}: color_data = 12'hd90;
			{8'd116, 8'd6}: color_data = 12'hd90;
			{8'd116, 8'd7}: color_data = 12'hea1;
			{8'd116, 8'd8}: color_data = 12'hfb4;
			{8'd116, 8'd9}: color_data = 12'hfc4;
			{8'd116, 8'd10}: color_data = 12'hea0;
			{8'd116, 8'd11}: color_data = 12'hd90;
			{8'd116, 8'd12}: color_data = 12'hd90;
			{8'd116, 8'd13}: color_data = 12'hd90;
			{8'd116, 8'd14}: color_data = 12'hd90;
			{8'd116, 8'd15}: color_data = 12'hea2;
			{8'd116, 8'd16}: color_data = 12'hfc5;
			{8'd116, 8'd17}: color_data = 12'hfc5;
			{8'd116, 8'd18}: color_data = 12'hfd5;
			{8'd116, 8'd55}: color_data = 12'h000;
			{8'd116, 8'd56}: color_data = 12'h763;
			{8'd116, 8'd57}: color_data = 12'hca5;
			{8'd116, 8'd58}: color_data = 12'h873;
			{8'd116, 8'd59}: color_data = 12'hfe7;
			{8'd116, 8'd60}: color_data = 12'hb95;
			{8'd116, 8'd61}: color_data = 12'hca8;
			{8'd116, 8'd62}: color_data = 12'hfdb;
			{8'd116, 8'd63}: color_data = 12'hfda;
			{8'd116, 8'd64}: color_data = 12'hfda;
			{8'd116, 8'd65}: color_data = 12'hfda;
			{8'd116, 8'd66}: color_data = 12'hfda;
			{8'd116, 8'd67}: color_data = 12'hfda;
			{8'd116, 8'd68}: color_data = 12'hfdb;
			{8'd116, 8'd69}: color_data = 12'hdb9;
			{8'd116, 8'd70}: color_data = 12'h865;
			{8'd116, 8'd71}: color_data = 12'hc97;
			{8'd116, 8'd72}: color_data = 12'hc97;
			{8'd116, 8'd73}: color_data = 12'hc97;
			{8'd116, 8'd74}: color_data = 12'hc97;
			{8'd116, 8'd75}: color_data = 12'hc97;
			{8'd116, 8'd76}: color_data = 12'h433;
			{8'd116, 8'd77}: color_data = 12'h012;
			{8'd116, 8'd78}: color_data = 12'h333;
			{8'd116, 8'd79}: color_data = 12'h865;
			{8'd116, 8'd80}: color_data = 12'hc97;
			{8'd116, 8'd81}: color_data = 12'hc97;
			{8'd116, 8'd82}: color_data = 12'hc97;
			{8'd116, 8'd83}: color_data = 12'hc97;
			{8'd116, 8'd84}: color_data = 12'hc97;
			{8'd116, 8'd85}: color_data = 12'hc97;
			{8'd116, 8'd86}: color_data = 12'hc97;
			{8'd116, 8'd87}: color_data = 12'hc97;
			{8'd116, 8'd88}: color_data = 12'hc97;
			{8'd116, 8'd89}: color_data = 12'hb97;
			{8'd116, 8'd90}: color_data = 12'h822;
			{8'd116, 8'd91}: color_data = 12'hf12;
			{8'd116, 8'd92}: color_data = 12'he12;
			{8'd116, 8'd93}: color_data = 12'he12;
			{8'd116, 8'd94}: color_data = 12'he12;
			{8'd116, 8'd95}: color_data = 12'he12;
			{8'd116, 8'd96}: color_data = 12'he12;
			{8'd116, 8'd97}: color_data = 12'he12;
			{8'd116, 8'd98}: color_data = 12'he12;
			{8'd116, 8'd99}: color_data = 12'hf12;
			{8'd116, 8'd100}: color_data = 12'ha11;
			{8'd116, 8'd101}: color_data = 12'h975;
			{8'd116, 8'd102}: color_data = 12'hc97;
			{8'd116, 8'd103}: color_data = 12'hc97;
			{8'd116, 8'd104}: color_data = 12'hc97;
			{8'd116, 8'd105}: color_data = 12'hc97;
			{8'd116, 8'd106}: color_data = 12'hc97;
			{8'd116, 8'd107}: color_data = 12'hc97;
			{8'd116, 8'd108}: color_data = 12'hc97;
			{8'd116, 8'd109}: color_data = 12'hc97;
			{8'd116, 8'd110}: color_data = 12'hc97;
			{8'd116, 8'd111}: color_data = 12'hc97;
			{8'd116, 8'd112}: color_data = 12'hc97;
			{8'd116, 8'd113}: color_data = 12'hc97;
			{8'd116, 8'd114}: color_data = 12'hc97;
			{8'd116, 8'd115}: color_data = 12'hc97;
			{8'd116, 8'd116}: color_data = 12'hc97;
			{8'd116, 8'd117}: color_data = 12'hc97;
			{8'd116, 8'd118}: color_data = 12'hc97;
			{8'd116, 8'd119}: color_data = 12'hc97;
			{8'd116, 8'd120}: color_data = 12'hc97;
			{8'd116, 8'd121}: color_data = 12'hc97;
			{8'd116, 8'd122}: color_data = 12'hc97;
			{8'd116, 8'd123}: color_data = 12'hc97;
			{8'd116, 8'd124}: color_data = 12'hc97;
			{8'd116, 8'd125}: color_data = 12'hc97;
			{8'd116, 8'd126}: color_data = 12'hc97;
			{8'd116, 8'd127}: color_data = 12'hd97;
			{8'd116, 8'd128}: color_data = 12'h754;
			{8'd116, 8'd129}: color_data = 12'h000;
			{8'd117, 8'd0}: color_data = 12'hfc4;
			{8'd117, 8'd1}: color_data = 12'hfc5;
			{8'd117, 8'd2}: color_data = 12'heb2;
			{8'd117, 8'd3}: color_data = 12'hd90;
			{8'd117, 8'd4}: color_data = 12'hd90;
			{8'd117, 8'd5}: color_data = 12'hd90;
			{8'd117, 8'd6}: color_data = 12'hd90;
			{8'd117, 8'd7}: color_data = 12'heb2;
			{8'd117, 8'd8}: color_data = 12'hfc5;
			{8'd117, 8'd9}: color_data = 12'hfc5;
			{8'd117, 8'd10}: color_data = 12'heb2;
			{8'd117, 8'd11}: color_data = 12'hd90;
			{8'd117, 8'd12}: color_data = 12'hd90;
			{8'd117, 8'd13}: color_data = 12'hd90;
			{8'd117, 8'd14}: color_data = 12'hd90;
			{8'd117, 8'd15}: color_data = 12'hd90;
			{8'd117, 8'd16}: color_data = 12'hfc4;
			{8'd117, 8'd17}: color_data = 12'hfc5;
			{8'd117, 8'd18}: color_data = 12'hfc5;
			{8'd117, 8'd55}: color_data = 12'h442;
			{8'd117, 8'd56}: color_data = 12'hb94;
			{8'd117, 8'd57}: color_data = 12'h763;
			{8'd117, 8'd58}: color_data = 12'hfd6;
			{8'd117, 8'd59}: color_data = 12'hfd6;
			{8'd117, 8'd60}: color_data = 12'hfd6;
			{8'd117, 8'd61}: color_data = 12'h984;
			{8'd117, 8'd62}: color_data = 12'hda9;
			{8'd117, 8'd63}: color_data = 12'hfdb;
			{8'd117, 8'd64}: color_data = 12'hfdb;
			{8'd117, 8'd65}: color_data = 12'hfdb;
			{8'd117, 8'd66}: color_data = 12'hfdb;
			{8'd117, 8'd67}: color_data = 12'hfca;
			{8'd117, 8'd68}: color_data = 12'hca8;
			{8'd117, 8'd69}: color_data = 12'h865;
			{8'd117, 8'd70}: color_data = 12'hb87;
			{8'd117, 8'd71}: color_data = 12'hc97;
			{8'd117, 8'd72}: color_data = 12'hc97;
			{8'd117, 8'd73}: color_data = 12'hc97;
			{8'd117, 8'd74}: color_data = 12'hc97;
			{8'd117, 8'd75}: color_data = 12'hb86;
			{8'd117, 8'd76}: color_data = 12'h223;
			{8'd117, 8'd77}: color_data = 12'h012;
			{8'd117, 8'd78}: color_data = 12'h755;
			{8'd117, 8'd79}: color_data = 12'ha86;
			{8'd117, 8'd80}: color_data = 12'h754;
			{8'd117, 8'd81}: color_data = 12'hb87;
			{8'd117, 8'd82}: color_data = 12'hc97;
			{8'd117, 8'd83}: color_data = 12'hc97;
			{8'd117, 8'd84}: color_data = 12'hc97;
			{8'd117, 8'd85}: color_data = 12'hc97;
			{8'd117, 8'd86}: color_data = 12'hc97;
			{8'd117, 8'd87}: color_data = 12'hc97;
			{8'd117, 8'd88}: color_data = 12'hc97;
			{8'd117, 8'd89}: color_data = 12'hc97;
			{8'd117, 8'd90}: color_data = 12'h975;
			{8'd117, 8'd91}: color_data = 12'ha11;
			{8'd117, 8'd92}: color_data = 12'hf12;
			{8'd117, 8'd93}: color_data = 12'hf12;
			{8'd117, 8'd94}: color_data = 12'he12;
			{8'd117, 8'd95}: color_data = 12'he12;
			{8'd117, 8'd96}: color_data = 12'he12;
			{8'd117, 8'd97}: color_data = 12'hf12;
			{8'd117, 8'd98}: color_data = 12'hf12;
			{8'd117, 8'd99}: color_data = 12'ha11;
			{8'd117, 8'd100}: color_data = 12'h854;
			{8'd117, 8'd101}: color_data = 12'hc97;
			{8'd117, 8'd102}: color_data = 12'hc97;
			{8'd117, 8'd103}: color_data = 12'hc97;
			{8'd117, 8'd104}: color_data = 12'hc97;
			{8'd117, 8'd105}: color_data = 12'hc97;
			{8'd117, 8'd106}: color_data = 12'hc97;
			{8'd117, 8'd107}: color_data = 12'hc97;
			{8'd117, 8'd108}: color_data = 12'hc97;
			{8'd117, 8'd109}: color_data = 12'hc97;
			{8'd117, 8'd110}: color_data = 12'hc97;
			{8'd117, 8'd111}: color_data = 12'hc97;
			{8'd117, 8'd112}: color_data = 12'hc97;
			{8'd117, 8'd113}: color_data = 12'hc97;
			{8'd117, 8'd114}: color_data = 12'hc97;
			{8'd117, 8'd115}: color_data = 12'hc97;
			{8'd117, 8'd116}: color_data = 12'hc97;
			{8'd117, 8'd117}: color_data = 12'hc97;
			{8'd117, 8'd118}: color_data = 12'hc97;
			{8'd117, 8'd119}: color_data = 12'hc97;
			{8'd117, 8'd120}: color_data = 12'hc97;
			{8'd117, 8'd121}: color_data = 12'hc97;
			{8'd117, 8'd122}: color_data = 12'hc97;
			{8'd117, 8'd123}: color_data = 12'hc97;
			{8'd117, 8'd124}: color_data = 12'hc97;
			{8'd117, 8'd125}: color_data = 12'hc97;
			{8'd117, 8'd126}: color_data = 12'hc97;
			{8'd117, 8'd127}: color_data = 12'hd97;
			{8'd117, 8'd128}: color_data = 12'h654;
			{8'd118, 8'd0}: color_data = 12'hfc5;
			{8'd118, 8'd1}: color_data = 12'hfc5;
			{8'd118, 8'd2}: color_data = 12'hea1;
			{8'd118, 8'd3}: color_data = 12'hd90;
			{8'd118, 8'd4}: color_data = 12'hd90;
			{8'd118, 8'd5}: color_data = 12'hd90;
			{8'd118, 8'd6}: color_data = 12'hd90;
			{8'd118, 8'd7}: color_data = 12'heb2;
			{8'd118, 8'd8}: color_data = 12'hfc6;
			{8'd118, 8'd9}: color_data = 12'hfc5;
			{8'd118, 8'd10}: color_data = 12'hea1;
			{8'd118, 8'd11}: color_data = 12'hd90;
			{8'd118, 8'd12}: color_data = 12'hd90;
			{8'd118, 8'd13}: color_data = 12'hd90;
			{8'd118, 8'd14}: color_data = 12'hd90;
			{8'd118, 8'd15}: color_data = 12'hd90;
			{8'd118, 8'd16}: color_data = 12'hfc5;
			{8'd118, 8'd17}: color_data = 12'hfc5;
			{8'd118, 8'd18}: color_data = 12'hfc5;
			{8'd118, 8'd55}: color_data = 12'h431;
			{8'd118, 8'd56}: color_data = 12'hb95;
			{8'd118, 8'd57}: color_data = 12'hca5;
			{8'd118, 8'd58}: color_data = 12'hfd7;
			{8'd118, 8'd59}: color_data = 12'hfd6;
			{8'd118, 8'd60}: color_data = 12'hfd6;
			{8'd118, 8'd61}: color_data = 12'hfd6;
			{8'd118, 8'd62}: color_data = 12'h984;
			{8'd118, 8'd63}: color_data = 12'h865;
			{8'd118, 8'd64}: color_data = 12'h986;
			{8'd118, 8'd65}: color_data = 12'hb97;
			{8'd118, 8'd66}: color_data = 12'h976;
			{8'd118, 8'd67}: color_data = 12'h875;
			{8'd118, 8'd68}: color_data = 12'h975;
			{8'd118, 8'd69}: color_data = 12'hc97;
			{8'd118, 8'd70}: color_data = 12'hc97;
			{8'd118, 8'd71}: color_data = 12'hc97;
			{8'd118, 8'd72}: color_data = 12'hc97;
			{8'd118, 8'd73}: color_data = 12'hc97;
			{8'd118, 8'd74}: color_data = 12'hc97;
			{8'd118, 8'd75}: color_data = 12'h975;
			{8'd118, 8'd76}: color_data = 12'h123;
			{8'd118, 8'd77}: color_data = 12'h112;
			{8'd118, 8'd78}: color_data = 12'h543;
			{8'd118, 8'd79}: color_data = 12'hc97;
			{8'd118, 8'd80}: color_data = 12'hb86;
			{8'd118, 8'd81}: color_data = 12'h754;
			{8'd118, 8'd82}: color_data = 12'h975;
			{8'd118, 8'd83}: color_data = 12'hc97;
			{8'd118, 8'd84}: color_data = 12'hc97;
			{8'd118, 8'd85}: color_data = 12'hc97;
			{8'd118, 8'd86}: color_data = 12'hc97;
			{8'd118, 8'd87}: color_data = 12'hc97;
			{8'd118, 8'd88}: color_data = 12'hc97;
			{8'd118, 8'd89}: color_data = 12'hc97;
			{8'd118, 8'd90}: color_data = 12'hc97;
			{8'd118, 8'd91}: color_data = 12'h965;
			{8'd118, 8'd92}: color_data = 12'h911;
			{8'd118, 8'd93}: color_data = 12'hd11;
			{8'd118, 8'd94}: color_data = 12'he12;
			{8'd118, 8'd95}: color_data = 12'he12;
			{8'd118, 8'd96}: color_data = 12'he11;
			{8'd118, 8'd97}: color_data = 12'hb11;
			{8'd118, 8'd98}: color_data = 12'h822;
			{8'd118, 8'd99}: color_data = 12'h975;
			{8'd118, 8'd100}: color_data = 12'hc97;
			{8'd118, 8'd101}: color_data = 12'hc97;
			{8'd118, 8'd102}: color_data = 12'hc97;
			{8'd118, 8'd103}: color_data = 12'hc97;
			{8'd118, 8'd104}: color_data = 12'hc97;
			{8'd118, 8'd105}: color_data = 12'hc97;
			{8'd118, 8'd106}: color_data = 12'hc97;
			{8'd118, 8'd107}: color_data = 12'hc97;
			{8'd118, 8'd108}: color_data = 12'hc97;
			{8'd118, 8'd109}: color_data = 12'hc97;
			{8'd118, 8'd110}: color_data = 12'hc97;
			{8'd118, 8'd111}: color_data = 12'hc97;
			{8'd118, 8'd112}: color_data = 12'hc97;
			{8'd118, 8'd113}: color_data = 12'hc97;
			{8'd118, 8'd114}: color_data = 12'hc97;
			{8'd118, 8'd115}: color_data = 12'hc97;
			{8'd118, 8'd116}: color_data = 12'hc97;
			{8'd118, 8'd117}: color_data = 12'hc97;
			{8'd118, 8'd118}: color_data = 12'hc97;
			{8'd118, 8'd119}: color_data = 12'hc97;
			{8'd118, 8'd120}: color_data = 12'hc97;
			{8'd118, 8'd121}: color_data = 12'hc97;
			{8'd118, 8'd122}: color_data = 12'hc97;
			{8'd118, 8'd123}: color_data = 12'ha76;
			{8'd118, 8'd124}: color_data = 12'hc97;
			{8'd118, 8'd125}: color_data = 12'hc97;
			{8'd118, 8'd126}: color_data = 12'hc97;
			{8'd118, 8'd127}: color_data = 12'hc97;
			{8'd118, 8'd128}: color_data = 12'h543;
			{8'd119, 8'd0}: color_data = 12'hfc5;
			{8'd119, 8'd1}: color_data = 12'hfc5;
			{8'd119, 8'd2}: color_data = 12'hea1;
			{8'd119, 8'd3}: color_data = 12'hd90;
			{8'd119, 8'd4}: color_data = 12'hd90;
			{8'd119, 8'd5}: color_data = 12'hd90;
			{8'd119, 8'd6}: color_data = 12'hd90;
			{8'd119, 8'd7}: color_data = 12'hd90;
			{8'd119, 8'd8}: color_data = 12'hea1;
			{8'd119, 8'd9}: color_data = 12'hea1;
			{8'd119, 8'd10}: color_data = 12'hd90;
			{8'd119, 8'd11}: color_data = 12'hd90;
			{8'd119, 8'd12}: color_data = 12'hd90;
			{8'd119, 8'd13}: color_data = 12'hd90;
			{8'd119, 8'd14}: color_data = 12'hd90;
			{8'd119, 8'd15}: color_data = 12'heb2;
			{8'd119, 8'd16}: color_data = 12'hfc5;
			{8'd119, 8'd17}: color_data = 12'hfc5;
			{8'd119, 8'd18}: color_data = 12'hfb4;
			{8'd119, 8'd55}: color_data = 12'h000;
			{8'd119, 8'd56}: color_data = 12'h431;
			{8'd119, 8'd57}: color_data = 12'hdc6;
			{8'd119, 8'd58}: color_data = 12'hfe7;
			{8'd119, 8'd59}: color_data = 12'hfe7;
			{8'd119, 8'd60}: color_data = 12'hfd6;
			{8'd119, 8'd61}: color_data = 12'hec6;
			{8'd119, 8'd62}: color_data = 12'h984;
			{8'd119, 8'd63}: color_data = 12'ha84;
			{8'd119, 8'd64}: color_data = 12'h652;
			{8'd119, 8'd65}: color_data = 12'hb94;
			{8'd119, 8'd66}: color_data = 12'h864;
			{8'd119, 8'd67}: color_data = 12'hc97;
			{8'd119, 8'd68}: color_data = 12'hc97;
			{8'd119, 8'd69}: color_data = 12'hc97;
			{8'd119, 8'd70}: color_data = 12'hc97;
			{8'd119, 8'd71}: color_data = 12'hc97;
			{8'd119, 8'd72}: color_data = 12'hc97;
			{8'd119, 8'd73}: color_data = 12'hc97;
			{8'd119, 8'd74}: color_data = 12'hd97;
			{8'd119, 8'd75}: color_data = 12'h754;
			{8'd119, 8'd76}: color_data = 12'h113;
			{8'd119, 8'd77}: color_data = 12'h222;
			{8'd119, 8'd78}: color_data = 12'h975;
			{8'd119, 8'd79}: color_data = 12'h865;
			{8'd119, 8'd80}: color_data = 12'hc97;
			{8'd119, 8'd81}: color_data = 12'hc97;
			{8'd119, 8'd82}: color_data = 12'h975;
			{8'd119, 8'd83}: color_data = 12'h764;
			{8'd119, 8'd84}: color_data = 12'h965;
			{8'd119, 8'd85}: color_data = 12'hc97;
			{8'd119, 8'd86}: color_data = 12'hc97;
			{8'd119, 8'd87}: color_data = 12'hc97;
			{8'd119, 8'd88}: color_data = 12'hc97;
			{8'd119, 8'd89}: color_data = 12'hc97;
			{8'd119, 8'd90}: color_data = 12'hc97;
			{8'd119, 8'd91}: color_data = 12'hc97;
			{8'd119, 8'd92}: color_data = 12'ha86;
			{8'd119, 8'd93}: color_data = 12'h854;
			{8'd119, 8'd94}: color_data = 12'h833;
			{8'd119, 8'd95}: color_data = 12'h833;
			{8'd119, 8'd96}: color_data = 12'h844;
			{8'd119, 8'd97}: color_data = 12'h975;
			{8'd119, 8'd98}: color_data = 12'hb97;
			{8'd119, 8'd99}: color_data = 12'hc97;
			{8'd119, 8'd100}: color_data = 12'hc97;
			{8'd119, 8'd101}: color_data = 12'hc97;
			{8'd119, 8'd102}: color_data = 12'hc97;
			{8'd119, 8'd103}: color_data = 12'hc97;
			{8'd119, 8'd104}: color_data = 12'hc97;
			{8'd119, 8'd105}: color_data = 12'hc97;
			{8'd119, 8'd106}: color_data = 12'hc97;
			{8'd119, 8'd107}: color_data = 12'hc97;
			{8'd119, 8'd108}: color_data = 12'hc97;
			{8'd119, 8'd109}: color_data = 12'hc97;
			{8'd119, 8'd110}: color_data = 12'hc97;
			{8'd119, 8'd111}: color_data = 12'hc97;
			{8'd119, 8'd112}: color_data = 12'hc97;
			{8'd119, 8'd113}: color_data = 12'hc97;
			{8'd119, 8'd114}: color_data = 12'hc97;
			{8'd119, 8'd115}: color_data = 12'hc97;
			{8'd119, 8'd116}: color_data = 12'hc97;
			{8'd119, 8'd117}: color_data = 12'hc97;
			{8'd119, 8'd118}: color_data = 12'hc97;
			{8'd119, 8'd119}: color_data = 12'hc97;
			{8'd119, 8'd120}: color_data = 12'hc97;
			{8'd119, 8'd121}: color_data = 12'hc97;
			{8'd119, 8'd122}: color_data = 12'hc97;
			{8'd119, 8'd123}: color_data = 12'h865;
			{8'd119, 8'd124}: color_data = 12'ha86;
			{8'd119, 8'd125}: color_data = 12'hc97;
			{8'd119, 8'd126}: color_data = 12'hc97;
			{8'd119, 8'd127}: color_data = 12'hc97;
			{8'd119, 8'd128}: color_data = 12'h322;
			{8'd120, 8'd0}: color_data = 12'hfc5;
			{8'd120, 8'd1}: color_data = 12'hfc5;
			{8'd120, 8'd2}: color_data = 12'hfc4;
			{8'd120, 8'd3}: color_data = 12'hda0;
			{8'd120, 8'd4}: color_data = 12'hd90;
			{8'd120, 8'd5}: color_data = 12'hd90;
			{8'd120, 8'd6}: color_data = 12'hd90;
			{8'd120, 8'd7}: color_data = 12'hd90;
			{8'd120, 8'd8}: color_data = 12'hd90;
			{8'd120, 8'd9}: color_data = 12'hd90;
			{8'd120, 8'd10}: color_data = 12'hd90;
			{8'd120, 8'd11}: color_data = 12'hd90;
			{8'd120, 8'd12}: color_data = 12'hd90;
			{8'd120, 8'd13}: color_data = 12'hd90;
			{8'd120, 8'd14}: color_data = 12'hd90;
			{8'd120, 8'd15}: color_data = 12'hfc4;
			{8'd120, 8'd16}: color_data = 12'hfc5;
			{8'd120, 8'd17}: color_data = 12'hfc5;
			{8'd120, 8'd56}: color_data = 12'h000;
			{8'd120, 8'd57}: color_data = 12'h763;
			{8'd120, 8'd58}: color_data = 12'hca5;
			{8'd120, 8'd59}: color_data = 12'hb94;
			{8'd120, 8'd60}: color_data = 12'ha84;
			{8'd120, 8'd61}: color_data = 12'ha94;
			{8'd120, 8'd62}: color_data = 12'h873;
			{8'd120, 8'd63}: color_data = 12'h873;
			{8'd120, 8'd64}: color_data = 12'hca5;
			{8'd120, 8'd65}: color_data = 12'h652;
			{8'd120, 8'd66}: color_data = 12'h754;
			{8'd120, 8'd67}: color_data = 12'hc97;
			{8'd120, 8'd68}: color_data = 12'hc97;
			{8'd120, 8'd69}: color_data = 12'hc97;
			{8'd120, 8'd70}: color_data = 12'hc97;
			{8'd120, 8'd71}: color_data = 12'hc97;
			{8'd120, 8'd72}: color_data = 12'hc97;
			{8'd120, 8'd73}: color_data = 12'hc97;
			{8'd120, 8'd74}: color_data = 12'hc97;
			{8'd120, 8'd75}: color_data = 12'h433;
			{8'd120, 8'd76}: color_data = 12'h113;
			{8'd120, 8'd77}: color_data = 12'h333;
			{8'd120, 8'd78}: color_data = 12'hc97;
			{8'd120, 8'd79}: color_data = 12'h965;
			{8'd120, 8'd80}: color_data = 12'h965;
			{8'd120, 8'd81}: color_data = 12'hd97;
			{8'd120, 8'd82}: color_data = 12'h975;
			{8'd120, 8'd83}: color_data = 12'ha86;
			{8'd120, 8'd84}: color_data = 12'hc97;
			{8'd120, 8'd85}: color_data = 12'hc97;
			{8'd120, 8'd86}: color_data = 12'hc97;
			{8'd120, 8'd87}: color_data = 12'hc97;
			{8'd120, 8'd88}: color_data = 12'hc97;
			{8'd120, 8'd89}: color_data = 12'hc97;
			{8'd120, 8'd90}: color_data = 12'hc97;
			{8'd120, 8'd91}: color_data = 12'hc97;
			{8'd120, 8'd92}: color_data = 12'hc97;
			{8'd120, 8'd93}: color_data = 12'hc97;
			{8'd120, 8'd94}: color_data = 12'hc97;
			{8'd120, 8'd95}: color_data = 12'hc97;
			{8'd120, 8'd96}: color_data = 12'hc97;
			{8'd120, 8'd97}: color_data = 12'hc97;
			{8'd120, 8'd98}: color_data = 12'hc97;
			{8'd120, 8'd99}: color_data = 12'hc97;
			{8'd120, 8'd100}: color_data = 12'hc97;
			{8'd120, 8'd101}: color_data = 12'hc97;
			{8'd120, 8'd102}: color_data = 12'hc97;
			{8'd120, 8'd103}: color_data = 12'hc97;
			{8'd120, 8'd104}: color_data = 12'hc97;
			{8'd120, 8'd105}: color_data = 12'hc97;
			{8'd120, 8'd106}: color_data = 12'hc97;
			{8'd120, 8'd107}: color_data = 12'hc97;
			{8'd120, 8'd108}: color_data = 12'hc97;
			{8'd120, 8'd109}: color_data = 12'hc97;
			{8'd120, 8'd110}: color_data = 12'hc97;
			{8'd120, 8'd111}: color_data = 12'hc97;
			{8'd120, 8'd112}: color_data = 12'hc97;
			{8'd120, 8'd113}: color_data = 12'hc97;
			{8'd120, 8'd114}: color_data = 12'hc97;
			{8'd120, 8'd115}: color_data = 12'hc97;
			{8'd120, 8'd116}: color_data = 12'hc97;
			{8'd120, 8'd117}: color_data = 12'hc97;
			{8'd120, 8'd118}: color_data = 12'hc97;
			{8'd120, 8'd119}: color_data = 12'hc97;
			{8'd120, 8'd120}: color_data = 12'hc97;
			{8'd120, 8'd121}: color_data = 12'hc97;
			{8'd120, 8'd122}: color_data = 12'hc97;
			{8'd120, 8'd123}: color_data = 12'ha76;
			{8'd120, 8'd124}: color_data = 12'h976;
			{8'd120, 8'd125}: color_data = 12'hc97;
			{8'd120, 8'd126}: color_data = 12'hc97;
			{8'd120, 8'd127}: color_data = 12'ha86;
			{8'd120, 8'd128}: color_data = 12'h110;
			{8'd121, 8'd0}: color_data = 12'hec4;
			{8'd121, 8'd1}: color_data = 12'hfc4;
			{8'd121, 8'd2}: color_data = 12'hfc5;
			{8'd121, 8'd3}: color_data = 12'hfb3;
			{8'd121, 8'd4}: color_data = 12'hd90;
			{8'd121, 8'd5}: color_data = 12'hd90;
			{8'd121, 8'd6}: color_data = 12'hd90;
			{8'd121, 8'd7}: color_data = 12'hd90;
			{8'd121, 8'd8}: color_data = 12'hd90;
			{8'd121, 8'd9}: color_data = 12'hd90;
			{8'd121, 8'd10}: color_data = 12'hd90;
			{8'd121, 8'd11}: color_data = 12'hd90;
			{8'd121, 8'd12}: color_data = 12'hd90;
			{8'd121, 8'd13}: color_data = 12'hd90;
			{8'd121, 8'd14}: color_data = 12'hea2;
			{8'd121, 8'd15}: color_data = 12'hfc5;
			{8'd121, 8'd16}: color_data = 12'hfc5;
			{8'd121, 8'd17}: color_data = 12'hfc6;
			{8'd121, 8'd57}: color_data = 12'h000;
			{8'd121, 8'd58}: color_data = 12'h000;
			{8'd121, 8'd59}: color_data = 12'h542;
			{8'd121, 8'd60}: color_data = 12'hfd6;
			{8'd121, 8'd61}: color_data = 12'hfd7;
			{8'd121, 8'd62}: color_data = 12'hfd6;
			{8'd121, 8'd63}: color_data = 12'h984;
			{8'd121, 8'd64}: color_data = 12'h763;
			{8'd121, 8'd65}: color_data = 12'h873;
			{8'd121, 8'd66}: color_data = 12'h653;
			{8'd121, 8'd67}: color_data = 12'hc97;
			{8'd121, 8'd68}: color_data = 12'hc97;
			{8'd121, 8'd69}: color_data = 12'hc97;
			{8'd121, 8'd70}: color_data = 12'hc97;
			{8'd121, 8'd71}: color_data = 12'hc97;
			{8'd121, 8'd72}: color_data = 12'hc97;
			{8'd121, 8'd73}: color_data = 12'hc97;
			{8'd121, 8'd74}: color_data = 12'h643;
			{8'd121, 8'd75}: color_data = 12'h001;
			{8'd121, 8'd76}: color_data = 12'h112;
			{8'd121, 8'd77}: color_data = 12'h544;
			{8'd121, 8'd78}: color_data = 12'hd97;
			{8'd121, 8'd79}: color_data = 12'hc97;
			{8'd121, 8'd80}: color_data = 12'h865;
			{8'd121, 8'd81}: color_data = 12'h975;
			{8'd121, 8'd82}: color_data = 12'hc97;
			{8'd121, 8'd83}: color_data = 12'h754;
			{8'd121, 8'd84}: color_data = 12'ha76;
			{8'd121, 8'd85}: color_data = 12'hc97;
			{8'd121, 8'd86}: color_data = 12'hc97;
			{8'd121, 8'd87}: color_data = 12'hc97;
			{8'd121, 8'd88}: color_data = 12'hc97;
			{8'd121, 8'd89}: color_data = 12'hc97;
			{8'd121, 8'd90}: color_data = 12'hc97;
			{8'd121, 8'd91}: color_data = 12'hc97;
			{8'd121, 8'd92}: color_data = 12'hc97;
			{8'd121, 8'd93}: color_data = 12'hc97;
			{8'd121, 8'd94}: color_data = 12'hc97;
			{8'd121, 8'd95}: color_data = 12'hc97;
			{8'd121, 8'd96}: color_data = 12'hc97;
			{8'd121, 8'd97}: color_data = 12'hc97;
			{8'd121, 8'd98}: color_data = 12'hc97;
			{8'd121, 8'd99}: color_data = 12'hc97;
			{8'd121, 8'd100}: color_data = 12'hc97;
			{8'd121, 8'd101}: color_data = 12'hc97;
			{8'd121, 8'd102}: color_data = 12'hc97;
			{8'd121, 8'd103}: color_data = 12'hc97;
			{8'd121, 8'd104}: color_data = 12'hc97;
			{8'd121, 8'd105}: color_data = 12'hc97;
			{8'd121, 8'd106}: color_data = 12'hc97;
			{8'd121, 8'd107}: color_data = 12'hc97;
			{8'd121, 8'd108}: color_data = 12'hc97;
			{8'd121, 8'd109}: color_data = 12'hc97;
			{8'd121, 8'd110}: color_data = 12'hc97;
			{8'd121, 8'd111}: color_data = 12'hc97;
			{8'd121, 8'd112}: color_data = 12'hc97;
			{8'd121, 8'd113}: color_data = 12'hc97;
			{8'd121, 8'd114}: color_data = 12'hc97;
			{8'd121, 8'd115}: color_data = 12'hc97;
			{8'd121, 8'd116}: color_data = 12'hc97;
			{8'd121, 8'd117}: color_data = 12'hc97;
			{8'd121, 8'd118}: color_data = 12'hc97;
			{8'd121, 8'd119}: color_data = 12'hc97;
			{8'd121, 8'd120}: color_data = 12'hc97;
			{8'd121, 8'd121}: color_data = 12'hc97;
			{8'd121, 8'd122}: color_data = 12'hc97;
			{8'd121, 8'd123}: color_data = 12'h865;
			{8'd121, 8'd124}: color_data = 12'ha86;
			{8'd121, 8'd125}: color_data = 12'hc97;
			{8'd121, 8'd126}: color_data = 12'hd97;
			{8'd121, 8'd127}: color_data = 12'h865;
			{8'd121, 8'd128}: color_data = 12'h000;
			{8'd122, 8'd1}: color_data = 12'hfc5;
			{8'd122, 8'd2}: color_data = 12'hfc4;
			{8'd122, 8'd3}: color_data = 12'hfc5;
			{8'd122, 8'd4}: color_data = 12'heb3;
			{8'd122, 8'd5}: color_data = 12'hd90;
			{8'd122, 8'd6}: color_data = 12'hd90;
			{8'd122, 8'd7}: color_data = 12'hd90;
			{8'd122, 8'd8}: color_data = 12'hd90;
			{8'd122, 8'd9}: color_data = 12'hd90;
			{8'd122, 8'd10}: color_data = 12'hd90;
			{8'd122, 8'd11}: color_data = 12'hd90;
			{8'd122, 8'd12}: color_data = 12'hd90;
			{8'd122, 8'd13}: color_data = 12'hd90;
			{8'd122, 8'd14}: color_data = 12'hfc4;
			{8'd122, 8'd15}: color_data = 12'hfc5;
			{8'd122, 8'd16}: color_data = 12'hfc5;
			{8'd122, 8'd59}: color_data = 12'h763;
			{8'd122, 8'd60}: color_data = 12'hfe7;
			{8'd122, 8'd61}: color_data = 12'hfd6;
			{8'd122, 8'd62}: color_data = 12'hfd6;
			{8'd122, 8'd63}: color_data = 12'hfd6;
			{8'd122, 8'd64}: color_data = 12'hec6;
			{8'd122, 8'd65}: color_data = 12'h652;
			{8'd122, 8'd66}: color_data = 12'h322;
			{8'd122, 8'd67}: color_data = 12'hc97;
			{8'd122, 8'd68}: color_data = 12'hc97;
			{8'd122, 8'd69}: color_data = 12'hc97;
			{8'd122, 8'd70}: color_data = 12'hc97;
			{8'd122, 8'd71}: color_data = 12'hc97;
			{8'd122, 8'd72}: color_data = 12'hc97;
			{8'd122, 8'd73}: color_data = 12'h543;
			{8'd122, 8'd74}: color_data = 12'h000;
			{8'd122, 8'd75}: color_data = 12'h000;
			{8'd122, 8'd76}: color_data = 12'h000;
			{8'd122, 8'd77}: color_data = 12'h432;
			{8'd122, 8'd78}: color_data = 12'hc97;
			{8'd122, 8'd79}: color_data = 12'hc97;
			{8'd122, 8'd80}: color_data = 12'hc97;
			{8'd122, 8'd81}: color_data = 12'h865;
			{8'd122, 8'd82}: color_data = 12'h865;
			{8'd122, 8'd83}: color_data = 12'hc97;
			{8'd122, 8'd84}: color_data = 12'h865;
			{8'd122, 8'd85}: color_data = 12'h975;
			{8'd122, 8'd86}: color_data = 12'hc97;
			{8'd122, 8'd87}: color_data = 12'hc97;
			{8'd122, 8'd88}: color_data = 12'hc97;
			{8'd122, 8'd89}: color_data = 12'hc97;
			{8'd122, 8'd90}: color_data = 12'hc97;
			{8'd122, 8'd91}: color_data = 12'hc97;
			{8'd122, 8'd92}: color_data = 12'hc97;
			{8'd122, 8'd93}: color_data = 12'hc97;
			{8'd122, 8'd94}: color_data = 12'hc97;
			{8'd122, 8'd95}: color_data = 12'hc97;
			{8'd122, 8'd96}: color_data = 12'hc97;
			{8'd122, 8'd97}: color_data = 12'hc97;
			{8'd122, 8'd98}: color_data = 12'hc97;
			{8'd122, 8'd99}: color_data = 12'hc97;
			{8'd122, 8'd100}: color_data = 12'hc97;
			{8'd122, 8'd101}: color_data = 12'hc97;
			{8'd122, 8'd102}: color_data = 12'hc97;
			{8'd122, 8'd103}: color_data = 12'hc97;
			{8'd122, 8'd104}: color_data = 12'hc97;
			{8'd122, 8'd105}: color_data = 12'hc97;
			{8'd122, 8'd106}: color_data = 12'hc97;
			{8'd122, 8'd107}: color_data = 12'hc97;
			{8'd122, 8'd108}: color_data = 12'hc97;
			{8'd122, 8'd109}: color_data = 12'hc97;
			{8'd122, 8'd110}: color_data = 12'hc97;
			{8'd122, 8'd111}: color_data = 12'hc97;
			{8'd122, 8'd112}: color_data = 12'hc97;
			{8'd122, 8'd113}: color_data = 12'hc97;
			{8'd122, 8'd114}: color_data = 12'hc97;
			{8'd122, 8'd115}: color_data = 12'hc97;
			{8'd122, 8'd116}: color_data = 12'hc97;
			{8'd122, 8'd117}: color_data = 12'hb87;
			{8'd122, 8'd118}: color_data = 12'h754;
			{8'd122, 8'd119}: color_data = 12'hc97;
			{8'd122, 8'd120}: color_data = 12'hc97;
			{8'd122, 8'd121}: color_data = 12'hc97;
			{8'd122, 8'd122}: color_data = 12'hb87;
			{8'd122, 8'd123}: color_data = 12'h754;
			{8'd122, 8'd124}: color_data = 12'hc97;
			{8'd122, 8'd125}: color_data = 12'hc97;
			{8'd122, 8'd126}: color_data = 12'hc97;
			{8'd122, 8'd127}: color_data = 12'h643;
			{8'd123, 8'd2}: color_data = 12'hfc5;
			{8'd123, 8'd3}: color_data = 12'hfc4;
			{8'd123, 8'd4}: color_data = 12'hfc5;
			{8'd123, 8'd5}: color_data = 12'heb2;
			{8'd123, 8'd6}: color_data = 12'hd90;
			{8'd123, 8'd7}: color_data = 12'hd90;
			{8'd123, 8'd8}: color_data = 12'hd90;
			{8'd123, 8'd9}: color_data = 12'hd90;
			{8'd123, 8'd10}: color_data = 12'hd90;
			{8'd123, 8'd11}: color_data = 12'hd90;
			{8'd123, 8'd12}: color_data = 12'hd90;
			{8'd123, 8'd13}: color_data = 12'hea1;
			{8'd123, 8'd14}: color_data = 12'hfc5;
			{8'd123, 8'd15}: color_data = 12'hfc5;
			{8'd123, 8'd16}: color_data = 12'hfc6;
			{8'd123, 8'd59}: color_data = 12'h321;
			{8'd123, 8'd60}: color_data = 12'hdb5;
			{8'd123, 8'd61}: color_data = 12'hfe7;
			{8'd123, 8'd62}: color_data = 12'hfe7;
			{8'd123, 8'd63}: color_data = 12'hfe7;
			{8'd123, 8'd64}: color_data = 12'hba5;
			{8'd123, 8'd65}: color_data = 12'h331;
			{8'd123, 8'd66}: color_data = 12'h000;
			{8'd123, 8'd67}: color_data = 12'ha76;
			{8'd123, 8'd68}: color_data = 12'hd97;
			{8'd123, 8'd69}: color_data = 12'hc97;
			{8'd123, 8'd70}: color_data = 12'hd97;
			{8'd123, 8'd71}: color_data = 12'hb86;
			{8'd123, 8'd72}: color_data = 12'h533;
			{8'd123, 8'd73}: color_data = 12'h000;
			{8'd123, 8'd77}: color_data = 12'h000;
			{8'd123, 8'd78}: color_data = 12'h754;
			{8'd123, 8'd79}: color_data = 12'hc97;
			{8'd123, 8'd80}: color_data = 12'hc97;
			{8'd123, 8'd81}: color_data = 12'hc97;
			{8'd123, 8'd82}: color_data = 12'ha76;
			{8'd123, 8'd83}: color_data = 12'h754;
			{8'd123, 8'd84}: color_data = 12'ha76;
			{8'd123, 8'd85}: color_data = 12'h865;
			{8'd123, 8'd86}: color_data = 12'ha76;
			{8'd123, 8'd87}: color_data = 12'hc97;
			{8'd123, 8'd88}: color_data = 12'hc97;
			{8'd123, 8'd89}: color_data = 12'hc97;
			{8'd123, 8'd90}: color_data = 12'hc97;
			{8'd123, 8'd91}: color_data = 12'hc97;
			{8'd123, 8'd92}: color_data = 12'hc97;
			{8'd123, 8'd93}: color_data = 12'hc97;
			{8'd123, 8'd94}: color_data = 12'hc97;
			{8'd123, 8'd95}: color_data = 12'hc97;
			{8'd123, 8'd96}: color_data = 12'hc97;
			{8'd123, 8'd97}: color_data = 12'hc97;
			{8'd123, 8'd98}: color_data = 12'hc97;
			{8'd123, 8'd99}: color_data = 12'hc97;
			{8'd123, 8'd100}: color_data = 12'hc97;
			{8'd123, 8'd101}: color_data = 12'hc97;
			{8'd123, 8'd102}: color_data = 12'hc97;
			{8'd123, 8'd103}: color_data = 12'hc97;
			{8'd123, 8'd104}: color_data = 12'hc97;
			{8'd123, 8'd105}: color_data = 12'hc97;
			{8'd123, 8'd106}: color_data = 12'hc97;
			{8'd123, 8'd107}: color_data = 12'hc97;
			{8'd123, 8'd108}: color_data = 12'hc97;
			{8'd123, 8'd109}: color_data = 12'hc97;
			{8'd123, 8'd110}: color_data = 12'hc97;
			{8'd123, 8'd111}: color_data = 12'hc97;
			{8'd123, 8'd112}: color_data = 12'hc97;
			{8'd123, 8'd113}: color_data = 12'hc97;
			{8'd123, 8'd114}: color_data = 12'hc97;
			{8'd123, 8'd115}: color_data = 12'hc97;
			{8'd123, 8'd116}: color_data = 12'hc97;
			{8'd123, 8'd117}: color_data = 12'h754;
			{8'd123, 8'd118}: color_data = 12'hb86;
			{8'd123, 8'd119}: color_data = 12'hc97;
			{8'd123, 8'd120}: color_data = 12'hc97;
			{8'd123, 8'd121}: color_data = 12'hc97;
			{8'd123, 8'd122}: color_data = 12'h764;
			{8'd123, 8'd123}: color_data = 12'hb86;
			{8'd123, 8'd124}: color_data = 12'hc97;
			{8'd123, 8'd125}: color_data = 12'hc97;
			{8'd123, 8'd126}: color_data = 12'hb86;
			{8'd123, 8'd127}: color_data = 12'h211;
			{8'd124, 8'd3}: color_data = 12'hfc5;
			{8'd124, 8'd4}: color_data = 12'hfc5;
			{8'd124, 8'd5}: color_data = 12'hfc5;
			{8'd124, 8'd6}: color_data = 12'hfb3;
			{8'd124, 8'd7}: color_data = 12'heb2;
			{8'd124, 8'd8}: color_data = 12'heb2;
			{8'd124, 8'd9}: color_data = 12'hea2;
			{8'd124, 8'd10}: color_data = 12'heb2;
			{8'd124, 8'd11}: color_data = 12'heb2;
			{8'd124, 8'd12}: color_data = 12'hea1;
			{8'd124, 8'd13}: color_data = 12'hfc4;
			{8'd124, 8'd14}: color_data = 12'hfc5;
			{8'd124, 8'd15}: color_data = 12'hfc5;
			{8'd124, 8'd59}: color_data = 12'h000;
			{8'd124, 8'd60}: color_data = 12'h321;
			{8'd124, 8'd61}: color_data = 12'h763;
			{8'd124, 8'd62}: color_data = 12'h973;
			{8'd124, 8'd63}: color_data = 12'h763;
			{8'd124, 8'd64}: color_data = 12'h210;
			{8'd124, 8'd66}: color_data = 12'h000;
			{8'd124, 8'd67}: color_data = 12'h432;
			{8'd124, 8'd68}: color_data = 12'h976;
			{8'd124, 8'd69}: color_data = 12'ha76;
			{8'd124, 8'd70}: color_data = 12'h754;
			{8'd124, 8'd71}: color_data = 12'h221;
			{8'd124, 8'd72}: color_data = 12'h000;
			{8'd124, 8'd78}: color_data = 12'h000;
			{8'd124, 8'd79}: color_data = 12'h865;
			{8'd124, 8'd80}: color_data = 12'hd97;
			{8'd124, 8'd81}: color_data = 12'hc97;
			{8'd124, 8'd82}: color_data = 12'hc97;
			{8'd124, 8'd83}: color_data = 12'hc97;
			{8'd124, 8'd84}: color_data = 12'h965;
			{8'd124, 8'd85}: color_data = 12'h754;
			{8'd124, 8'd86}: color_data = 12'h543;
			{8'd124, 8'd87}: color_data = 12'hb87;
			{8'd124, 8'd88}: color_data = 12'hc97;
			{8'd124, 8'd89}: color_data = 12'hc97;
			{8'd124, 8'd90}: color_data = 12'hc97;
			{8'd124, 8'd91}: color_data = 12'hc97;
			{8'd124, 8'd92}: color_data = 12'hc97;
			{8'd124, 8'd93}: color_data = 12'hc97;
			{8'd124, 8'd94}: color_data = 12'hc97;
			{8'd124, 8'd95}: color_data = 12'hc97;
			{8'd124, 8'd96}: color_data = 12'hc97;
			{8'd124, 8'd97}: color_data = 12'hc97;
			{8'd124, 8'd98}: color_data = 12'hc97;
			{8'd124, 8'd99}: color_data = 12'hc97;
			{8'd124, 8'd100}: color_data = 12'hc97;
			{8'd124, 8'd101}: color_data = 12'hc97;
			{8'd124, 8'd102}: color_data = 12'hc97;
			{8'd124, 8'd103}: color_data = 12'hc97;
			{8'd124, 8'd104}: color_data = 12'hc97;
			{8'd124, 8'd105}: color_data = 12'hc97;
			{8'd124, 8'd106}: color_data = 12'hc97;
			{8'd124, 8'd107}: color_data = 12'hc97;
			{8'd124, 8'd108}: color_data = 12'hc97;
			{8'd124, 8'd109}: color_data = 12'hc97;
			{8'd124, 8'd110}: color_data = 12'hc97;
			{8'd124, 8'd111}: color_data = 12'hc97;
			{8'd124, 8'd112}: color_data = 12'hc97;
			{8'd124, 8'd113}: color_data = 12'hc97;
			{8'd124, 8'd114}: color_data = 12'hc97;
			{8'd124, 8'd115}: color_data = 12'hb86;
			{8'd124, 8'd116}: color_data = 12'h754;
			{8'd124, 8'd117}: color_data = 12'hb86;
			{8'd124, 8'd118}: color_data = 12'hc97;
			{8'd124, 8'd119}: color_data = 12'hc97;
			{8'd124, 8'd120}: color_data = 12'hc97;
			{8'd124, 8'd121}: color_data = 12'h965;
			{8'd124, 8'd122}: color_data = 12'h975;
			{8'd124, 8'd123}: color_data = 12'hc97;
			{8'd124, 8'd124}: color_data = 12'hc97;
			{8'd124, 8'd125}: color_data = 12'hd97;
			{8'd124, 8'd126}: color_data = 12'h754;
			{8'd124, 8'd127}: color_data = 12'h000;
			{8'd125, 8'd4}: color_data = 12'hfc5;
			{8'd125, 8'd5}: color_data = 12'hfc5;
			{8'd125, 8'd6}: color_data = 12'hfc5;
			{8'd125, 8'd7}: color_data = 12'hfc5;
			{8'd125, 8'd8}: color_data = 12'hfc5;
			{8'd125, 8'd9}: color_data = 12'hfc5;
			{8'd125, 8'd10}: color_data = 12'hfc5;
			{8'd125, 8'd11}: color_data = 12'hfc6;
			{8'd125, 8'd12}: color_data = 12'hfc6;
			{8'd125, 8'd13}: color_data = 12'hfc5;
			{8'd125, 8'd14}: color_data = 12'hfc4;
			{8'd125, 8'd15}: color_data = 12'hfb3;
			{8'd125, 8'd62}: color_data = 12'h000;
			{8'd125, 8'd67}: color_data = 12'h000;
			{8'd125, 8'd68}: color_data = 12'h000;
			{8'd125, 8'd69}: color_data = 12'h000;
			{8'd125, 8'd70}: color_data = 12'h000;
			{8'd125, 8'd79}: color_data = 12'h111;
			{8'd125, 8'd80}: color_data = 12'h975;
			{8'd125, 8'd81}: color_data = 12'hd97;
			{8'd125, 8'd82}: color_data = 12'hc97;
			{8'd125, 8'd83}: color_data = 12'hc97;
			{8'd125, 8'd84}: color_data = 12'hc97;
			{8'd125, 8'd85}: color_data = 12'hc97;
			{8'd125, 8'd86}: color_data = 12'hb86;
			{8'd125, 8'd87}: color_data = 12'hc97;
			{8'd125, 8'd88}: color_data = 12'hc97;
			{8'd125, 8'd89}: color_data = 12'hc97;
			{8'd125, 8'd90}: color_data = 12'hc97;
			{8'd125, 8'd91}: color_data = 12'hc97;
			{8'd125, 8'd92}: color_data = 12'hc97;
			{8'd125, 8'd93}: color_data = 12'hc97;
			{8'd125, 8'd94}: color_data = 12'hc97;
			{8'd125, 8'd95}: color_data = 12'hc97;
			{8'd125, 8'd96}: color_data = 12'hc97;
			{8'd125, 8'd97}: color_data = 12'hc97;
			{8'd125, 8'd98}: color_data = 12'hc97;
			{8'd125, 8'd99}: color_data = 12'hc97;
			{8'd125, 8'd100}: color_data = 12'hc97;
			{8'd125, 8'd101}: color_data = 12'hc97;
			{8'd125, 8'd102}: color_data = 12'hc97;
			{8'd125, 8'd103}: color_data = 12'hc97;
			{8'd125, 8'd104}: color_data = 12'hc97;
			{8'd125, 8'd105}: color_data = 12'hc97;
			{8'd125, 8'd106}: color_data = 12'hc97;
			{8'd125, 8'd107}: color_data = 12'hc97;
			{8'd125, 8'd108}: color_data = 12'hc97;
			{8'd125, 8'd109}: color_data = 12'hc97;
			{8'd125, 8'd110}: color_data = 12'hc97;
			{8'd125, 8'd111}: color_data = 12'hc97;
			{8'd125, 8'd112}: color_data = 12'hc97;
			{8'd125, 8'd113}: color_data = 12'hb87;
			{8'd125, 8'd114}: color_data = 12'h975;
			{8'd125, 8'd115}: color_data = 12'h754;
			{8'd125, 8'd116}: color_data = 12'hb87;
			{8'd125, 8'd117}: color_data = 12'hc97;
			{8'd125, 8'd118}: color_data = 12'hc97;
			{8'd125, 8'd119}: color_data = 12'hc97;
			{8'd125, 8'd120}: color_data = 12'h976;
			{8'd125, 8'd121}: color_data = 12'h865;
			{8'd125, 8'd122}: color_data = 12'hc97;
			{8'd125, 8'd123}: color_data = 12'hc97;
			{8'd125, 8'd124}: color_data = 12'hc97;
			{8'd125, 8'd125}: color_data = 12'hb86;
			{8'd125, 8'd126}: color_data = 12'h321;
			{8'd126, 8'd5}: color_data = 12'hfc5;
			{8'd126, 8'd6}: color_data = 12'hfc5;
			{8'd126, 8'd7}: color_data = 12'hfc5;
			{8'd126, 8'd8}: color_data = 12'hfc5;
			{8'd126, 8'd9}: color_data = 12'hfc5;
			{8'd126, 8'd10}: color_data = 12'hfc5;
			{8'd126, 8'd11}: color_data = 12'hfc5;
			{8'd126, 8'd12}: color_data = 12'hfc5;
			{8'd126, 8'd13}: color_data = 12'hfc5;
			{8'd126, 8'd14}: color_data = 12'hfc5;
			{8'd126, 8'd80}: color_data = 12'h322;
			{8'd126, 8'd81}: color_data = 12'ha86;
			{8'd126, 8'd82}: color_data = 12'hc97;
			{8'd126, 8'd83}: color_data = 12'hc97;
			{8'd126, 8'd84}: color_data = 12'hc97;
			{8'd126, 8'd85}: color_data = 12'hc97;
			{8'd126, 8'd86}: color_data = 12'hc97;
			{8'd126, 8'd87}: color_data = 12'hc97;
			{8'd126, 8'd88}: color_data = 12'hc97;
			{8'd126, 8'd89}: color_data = 12'hc97;
			{8'd126, 8'd90}: color_data = 12'hc97;
			{8'd126, 8'd91}: color_data = 12'hc97;
			{8'd126, 8'd92}: color_data = 12'hc97;
			{8'd126, 8'd93}: color_data = 12'hc97;
			{8'd126, 8'd94}: color_data = 12'hc97;
			{8'd126, 8'd95}: color_data = 12'hc97;
			{8'd126, 8'd96}: color_data = 12'hc97;
			{8'd126, 8'd97}: color_data = 12'hc97;
			{8'd126, 8'd98}: color_data = 12'hc97;
			{8'd126, 8'd99}: color_data = 12'hc97;
			{8'd126, 8'd100}: color_data = 12'hc97;
			{8'd126, 8'd101}: color_data = 12'hc97;
			{8'd126, 8'd102}: color_data = 12'hc97;
			{8'd126, 8'd103}: color_data = 12'hc97;
			{8'd126, 8'd104}: color_data = 12'hc97;
			{8'd126, 8'd105}: color_data = 12'hc97;
			{8'd126, 8'd106}: color_data = 12'hc97;
			{8'd126, 8'd107}: color_data = 12'hc97;
			{8'd126, 8'd108}: color_data = 12'hc97;
			{8'd126, 8'd109}: color_data = 12'hc97;
			{8'd126, 8'd110}: color_data = 12'hc97;
			{8'd126, 8'd111}: color_data = 12'h965;
			{8'd126, 8'd112}: color_data = 12'h754;
			{8'd126, 8'd113}: color_data = 12'h864;
			{8'd126, 8'd114}: color_data = 12'ha76;
			{8'd126, 8'd115}: color_data = 12'hc97;
			{8'd126, 8'd116}: color_data = 12'hc97;
			{8'd126, 8'd117}: color_data = 12'hc97;
			{8'd126, 8'd118}: color_data = 12'hc97;
			{8'd126, 8'd119}: color_data = 12'h975;
			{8'd126, 8'd120}: color_data = 12'h864;
			{8'd126, 8'd121}: color_data = 12'hc97;
			{8'd126, 8'd122}: color_data = 12'hc97;
			{8'd126, 8'd123}: color_data = 12'hc97;
			{8'd126, 8'd124}: color_data = 12'hc97;
			{8'd126, 8'd125}: color_data = 12'h643;
			{8'd126, 8'd126}: color_data = 12'h000;
			{8'd127, 8'd81}: color_data = 12'h432;
			{8'd127, 8'd82}: color_data = 12'hb87;
			{8'd127, 8'd83}: color_data = 12'hc97;
			{8'd127, 8'd84}: color_data = 12'hc97;
			{8'd127, 8'd85}: color_data = 12'hc97;
			{8'd127, 8'd86}: color_data = 12'hc97;
			{8'd127, 8'd87}: color_data = 12'hc97;
			{8'd127, 8'd88}: color_data = 12'hc97;
			{8'd127, 8'd89}: color_data = 12'hc97;
			{8'd127, 8'd90}: color_data = 12'hc97;
			{8'd127, 8'd91}: color_data = 12'hc97;
			{8'd127, 8'd92}: color_data = 12'hc97;
			{8'd127, 8'd93}: color_data = 12'hc97;
			{8'd127, 8'd94}: color_data = 12'hc97;
			{8'd127, 8'd95}: color_data = 12'hc97;
			{8'd127, 8'd96}: color_data = 12'hc97;
			{8'd127, 8'd97}: color_data = 12'hc97;
			{8'd127, 8'd98}: color_data = 12'hc97;
			{8'd127, 8'd99}: color_data = 12'hc97;
			{8'd127, 8'd100}: color_data = 12'hc97;
			{8'd127, 8'd101}: color_data = 12'hc97;
			{8'd127, 8'd102}: color_data = 12'hc97;
			{8'd127, 8'd103}: color_data = 12'hc97;
			{8'd127, 8'd104}: color_data = 12'hc97;
			{8'd127, 8'd105}: color_data = 12'hc97;
			{8'd127, 8'd106}: color_data = 12'hc97;
			{8'd127, 8'd107}: color_data = 12'hc97;
			{8'd127, 8'd108}: color_data = 12'hc97;
			{8'd127, 8'd109}: color_data = 12'hc97;
			{8'd127, 8'd110}: color_data = 12'hc97;
			{8'd127, 8'd111}: color_data = 12'hb87;
			{8'd127, 8'd112}: color_data = 12'hc97;
			{8'd127, 8'd113}: color_data = 12'hc97;
			{8'd127, 8'd114}: color_data = 12'hc97;
			{8'd127, 8'd115}: color_data = 12'hc97;
			{8'd127, 8'd116}: color_data = 12'hc97;
			{8'd127, 8'd117}: color_data = 12'hc97;
			{8'd127, 8'd118}: color_data = 12'h865;
			{8'd127, 8'd119}: color_data = 12'h865;
			{8'd127, 8'd120}: color_data = 12'hc97;
			{8'd127, 8'd121}: color_data = 12'hc97;
			{8'd127, 8'd122}: color_data = 12'hc97;
			{8'd127, 8'd123}: color_data = 12'hd97;
			{8'd127, 8'd124}: color_data = 12'h865;
			{8'd127, 8'd125}: color_data = 12'h000;
			{8'd128, 8'd81}: color_data = 12'h000;
			{8'd128, 8'd82}: color_data = 12'h533;
			{8'd128, 8'd83}: color_data = 12'hc97;
			{8'd128, 8'd84}: color_data = 12'hc97;
			{8'd128, 8'd85}: color_data = 12'hc97;
			{8'd128, 8'd86}: color_data = 12'hc97;
			{8'd128, 8'd87}: color_data = 12'hc97;
			{8'd128, 8'd88}: color_data = 12'hc97;
			{8'd128, 8'd89}: color_data = 12'hc97;
			{8'd128, 8'd90}: color_data = 12'hc97;
			{8'd128, 8'd91}: color_data = 12'hc97;
			{8'd128, 8'd92}: color_data = 12'hc97;
			{8'd128, 8'd93}: color_data = 12'hc97;
			{8'd128, 8'd94}: color_data = 12'hc97;
			{8'd128, 8'd95}: color_data = 12'hc97;
			{8'd128, 8'd96}: color_data = 12'hc97;
			{8'd128, 8'd97}: color_data = 12'hc97;
			{8'd128, 8'd98}: color_data = 12'hc97;
			{8'd128, 8'd99}: color_data = 12'hc97;
			{8'd128, 8'd100}: color_data = 12'hc97;
			{8'd128, 8'd101}: color_data = 12'hc97;
			{8'd128, 8'd102}: color_data = 12'hc97;
			{8'd128, 8'd103}: color_data = 12'hc97;
			{8'd128, 8'd104}: color_data = 12'hc97;
			{8'd128, 8'd105}: color_data = 12'hc97;
			{8'd128, 8'd106}: color_data = 12'hc97;
			{8'd128, 8'd107}: color_data = 12'hc97;
			{8'd128, 8'd108}: color_data = 12'hc97;
			{8'd128, 8'd109}: color_data = 12'hc97;
			{8'd128, 8'd110}: color_data = 12'hc97;
			{8'd128, 8'd111}: color_data = 12'hc97;
			{8'd128, 8'd112}: color_data = 12'hc97;
			{8'd128, 8'd113}: color_data = 12'hc97;
			{8'd128, 8'd114}: color_data = 12'hc97;
			{8'd128, 8'd115}: color_data = 12'hc97;
			{8'd128, 8'd116}: color_data = 12'hc97;
			{8'd128, 8'd117}: color_data = 12'h864;
			{8'd128, 8'd118}: color_data = 12'h975;
			{8'd128, 8'd119}: color_data = 12'hc97;
			{8'd128, 8'd120}: color_data = 12'hc97;
			{8'd128, 8'd121}: color_data = 12'hc97;
			{8'd128, 8'd122}: color_data = 12'hd97;
			{8'd128, 8'd123}: color_data = 12'h975;
			{8'd128, 8'd124}: color_data = 12'h211;
			{8'd129, 8'd82}: color_data = 12'h000;
			{8'd129, 8'd83}: color_data = 12'h543;
			{8'd129, 8'd84}: color_data = 12'hc97;
			{8'd129, 8'd85}: color_data = 12'hc97;
			{8'd129, 8'd86}: color_data = 12'hc97;
			{8'd129, 8'd87}: color_data = 12'hc97;
			{8'd129, 8'd88}: color_data = 12'hc97;
			{8'd129, 8'd89}: color_data = 12'hc97;
			{8'd129, 8'd90}: color_data = 12'hc97;
			{8'd129, 8'd91}: color_data = 12'hc97;
			{8'd129, 8'd92}: color_data = 12'hc97;
			{8'd129, 8'd93}: color_data = 12'hc97;
			{8'd129, 8'd94}: color_data = 12'hc97;
			{8'd129, 8'd95}: color_data = 12'hc97;
			{8'd129, 8'd96}: color_data = 12'hc97;
			{8'd129, 8'd97}: color_data = 12'hc97;
			{8'd129, 8'd98}: color_data = 12'hc97;
			{8'd129, 8'd99}: color_data = 12'hc97;
			{8'd129, 8'd100}: color_data = 12'hc97;
			{8'd129, 8'd101}: color_data = 12'hc97;
			{8'd129, 8'd102}: color_data = 12'hc97;
			{8'd129, 8'd103}: color_data = 12'hc97;
			{8'd129, 8'd104}: color_data = 12'hc97;
			{8'd129, 8'd105}: color_data = 12'hc97;
			{8'd129, 8'd106}: color_data = 12'hc97;
			{8'd129, 8'd107}: color_data = 12'hc97;
			{8'd129, 8'd108}: color_data = 12'hc97;
			{8'd129, 8'd109}: color_data = 12'hc97;
			{8'd129, 8'd110}: color_data = 12'hc97;
			{8'd129, 8'd111}: color_data = 12'hc97;
			{8'd129, 8'd112}: color_data = 12'hc97;
			{8'd129, 8'd113}: color_data = 12'hc97;
			{8'd129, 8'd114}: color_data = 12'hc97;
			{8'd129, 8'd115}: color_data = 12'hc97;
			{8'd129, 8'd116}: color_data = 12'hc97;
			{8'd129, 8'd117}: color_data = 12'hb87;
			{8'd129, 8'd118}: color_data = 12'hc97;
			{8'd129, 8'd119}: color_data = 12'hc97;
			{8'd129, 8'd120}: color_data = 12'hc97;
			{8'd129, 8'd121}: color_data = 12'hd97;
			{8'd129, 8'd122}: color_data = 12'h975;
			{8'd129, 8'd123}: color_data = 12'h221;
			{8'd130, 8'd83}: color_data = 12'h000;
			{8'd130, 8'd84}: color_data = 12'h643;
			{8'd130, 8'd85}: color_data = 12'hc97;
			{8'd130, 8'd86}: color_data = 12'hc97;
			{8'd130, 8'd87}: color_data = 12'hc97;
			{8'd130, 8'd88}: color_data = 12'hc97;
			{8'd130, 8'd89}: color_data = 12'hc97;
			{8'd130, 8'd90}: color_data = 12'hc97;
			{8'd130, 8'd91}: color_data = 12'hc97;
			{8'd130, 8'd92}: color_data = 12'hc97;
			{8'd130, 8'd93}: color_data = 12'hc97;
			{8'd130, 8'd94}: color_data = 12'hc97;
			{8'd130, 8'd95}: color_data = 12'hc97;
			{8'd130, 8'd96}: color_data = 12'hc97;
			{8'd130, 8'd97}: color_data = 12'hc97;
			{8'd130, 8'd98}: color_data = 12'hc97;
			{8'd130, 8'd99}: color_data = 12'hc97;
			{8'd130, 8'd100}: color_data = 12'hc97;
			{8'd130, 8'd101}: color_data = 12'hc97;
			{8'd130, 8'd102}: color_data = 12'hc97;
			{8'd130, 8'd103}: color_data = 12'hc97;
			{8'd130, 8'd104}: color_data = 12'hc97;
			{8'd130, 8'd105}: color_data = 12'hc97;
			{8'd130, 8'd106}: color_data = 12'hc97;
			{8'd130, 8'd107}: color_data = 12'hc97;
			{8'd130, 8'd108}: color_data = 12'hc97;
			{8'd130, 8'd109}: color_data = 12'hc97;
			{8'd130, 8'd110}: color_data = 12'hc97;
			{8'd130, 8'd111}: color_data = 12'hc97;
			{8'd130, 8'd112}: color_data = 12'hc97;
			{8'd130, 8'd113}: color_data = 12'hc97;
			{8'd130, 8'd114}: color_data = 12'hc97;
			{8'd130, 8'd115}: color_data = 12'hc97;
			{8'd130, 8'd116}: color_data = 12'hc97;
			{8'd130, 8'd117}: color_data = 12'hc97;
			{8'd130, 8'd118}: color_data = 12'hc97;
			{8'd130, 8'd119}: color_data = 12'hc97;
			{8'd130, 8'd120}: color_data = 12'hd97;
			{8'd130, 8'd121}: color_data = 12'h865;
			{8'd130, 8'd122}: color_data = 12'h211;
			{8'd131, 8'd84}: color_data = 12'h000;
			{8'd131, 8'd85}: color_data = 12'h643;
			{8'd131, 8'd86}: color_data = 12'hc97;
			{8'd131, 8'd87}: color_data = 12'hc97;
			{8'd131, 8'd88}: color_data = 12'hc97;
			{8'd131, 8'd89}: color_data = 12'hc97;
			{8'd131, 8'd90}: color_data = 12'hc97;
			{8'd131, 8'd91}: color_data = 12'hc97;
			{8'd131, 8'd92}: color_data = 12'hc97;
			{8'd131, 8'd93}: color_data = 12'hc97;
			{8'd131, 8'd94}: color_data = 12'hc97;
			{8'd131, 8'd95}: color_data = 12'hc97;
			{8'd131, 8'd96}: color_data = 12'hc97;
			{8'd131, 8'd97}: color_data = 12'hc97;
			{8'd131, 8'd98}: color_data = 12'hc97;
			{8'd131, 8'd99}: color_data = 12'hc97;
			{8'd131, 8'd100}: color_data = 12'hc97;
			{8'd131, 8'd101}: color_data = 12'hc97;
			{8'd131, 8'd102}: color_data = 12'hc97;
			{8'd131, 8'd103}: color_data = 12'hc97;
			{8'd131, 8'd104}: color_data = 12'hc97;
			{8'd131, 8'd105}: color_data = 12'hc97;
			{8'd131, 8'd106}: color_data = 12'hc97;
			{8'd131, 8'd107}: color_data = 12'hc97;
			{8'd131, 8'd108}: color_data = 12'hc97;
			{8'd131, 8'd109}: color_data = 12'hc97;
			{8'd131, 8'd110}: color_data = 12'hc97;
			{8'd131, 8'd111}: color_data = 12'hc97;
			{8'd131, 8'd112}: color_data = 12'hc97;
			{8'd131, 8'd113}: color_data = 12'hc97;
			{8'd131, 8'd114}: color_data = 12'hc97;
			{8'd131, 8'd115}: color_data = 12'hc97;
			{8'd131, 8'd116}: color_data = 12'hc97;
			{8'd131, 8'd117}: color_data = 12'hc97;
			{8'd131, 8'd118}: color_data = 12'hc97;
			{8'd131, 8'd119}: color_data = 12'hc97;
			{8'd131, 8'd120}: color_data = 12'h754;
			{8'd131, 8'd121}: color_data = 12'h000;
			{8'd132, 8'd85}: color_data = 12'h000;
			{8'd132, 8'd86}: color_data = 12'h543;
			{8'd132, 8'd87}: color_data = 12'hb87;
			{8'd132, 8'd88}: color_data = 12'hc97;
			{8'd132, 8'd89}: color_data = 12'hc97;
			{8'd132, 8'd90}: color_data = 12'hc97;
			{8'd132, 8'd91}: color_data = 12'hc97;
			{8'd132, 8'd92}: color_data = 12'hc97;
			{8'd132, 8'd93}: color_data = 12'hc97;
			{8'd132, 8'd94}: color_data = 12'hc97;
			{8'd132, 8'd95}: color_data = 12'hc97;
			{8'd132, 8'd96}: color_data = 12'hc97;
			{8'd132, 8'd97}: color_data = 12'hc97;
			{8'd132, 8'd98}: color_data = 12'hc97;
			{8'd132, 8'd99}: color_data = 12'hc97;
			{8'd132, 8'd100}: color_data = 12'hc97;
			{8'd132, 8'd101}: color_data = 12'hc97;
			{8'd132, 8'd102}: color_data = 12'hc97;
			{8'd132, 8'd103}: color_data = 12'hc97;
			{8'd132, 8'd104}: color_data = 12'hc97;
			{8'd132, 8'd105}: color_data = 12'hc97;
			{8'd132, 8'd106}: color_data = 12'hc97;
			{8'd132, 8'd107}: color_data = 12'hc97;
			{8'd132, 8'd108}: color_data = 12'hc97;
			{8'd132, 8'd109}: color_data = 12'hc97;
			{8'd132, 8'd110}: color_data = 12'hc97;
			{8'd132, 8'd111}: color_data = 12'hc97;
			{8'd132, 8'd112}: color_data = 12'hc97;
			{8'd132, 8'd113}: color_data = 12'hc97;
			{8'd132, 8'd114}: color_data = 12'hc97;
			{8'd132, 8'd115}: color_data = 12'hc97;
			{8'd132, 8'd116}: color_data = 12'hc97;
			{8'd132, 8'd117}: color_data = 12'hd97;
			{8'd132, 8'd118}: color_data = 12'ha86;
			{8'd132, 8'd119}: color_data = 12'h533;
			{8'd132, 8'd120}: color_data = 12'h000;
			{8'd133, 8'd86}: color_data = 12'h000;
			{8'd133, 8'd87}: color_data = 12'h322;
			{8'd133, 8'd88}: color_data = 12'h975;
			{8'd133, 8'd89}: color_data = 12'hd97;
			{8'd133, 8'd90}: color_data = 12'hc97;
			{8'd133, 8'd91}: color_data = 12'hc97;
			{8'd133, 8'd92}: color_data = 12'hc97;
			{8'd133, 8'd93}: color_data = 12'hc97;
			{8'd133, 8'd94}: color_data = 12'hc97;
			{8'd133, 8'd95}: color_data = 12'hc97;
			{8'd133, 8'd96}: color_data = 12'hc97;
			{8'd133, 8'd97}: color_data = 12'hc97;
			{8'd133, 8'd98}: color_data = 12'hc97;
			{8'd133, 8'd99}: color_data = 12'hc97;
			{8'd133, 8'd100}: color_data = 12'hc97;
			{8'd133, 8'd101}: color_data = 12'hc97;
			{8'd133, 8'd102}: color_data = 12'hc97;
			{8'd133, 8'd103}: color_data = 12'hc97;
			{8'd133, 8'd104}: color_data = 12'hc97;
			{8'd133, 8'd105}: color_data = 12'hc97;
			{8'd133, 8'd106}: color_data = 12'hc97;
			{8'd133, 8'd107}: color_data = 12'hc97;
			{8'd133, 8'd108}: color_data = 12'hc97;
			{8'd133, 8'd109}: color_data = 12'hc97;
			{8'd133, 8'd110}: color_data = 12'hc97;
			{8'd133, 8'd111}: color_data = 12'hc97;
			{8'd133, 8'd112}: color_data = 12'hc97;
			{8'd133, 8'd113}: color_data = 12'hc97;
			{8'd133, 8'd114}: color_data = 12'hc97;
			{8'd133, 8'd115}: color_data = 12'hd97;
			{8'd133, 8'd116}: color_data = 12'hc97;
			{8'd133, 8'd117}: color_data = 12'h754;
			{8'd133, 8'd118}: color_data = 12'h211;
			{8'd133, 8'd119}: color_data = 12'h000;
			{8'd134, 8'd88}: color_data = 12'h100;
			{8'd134, 8'd89}: color_data = 12'h643;
			{8'd134, 8'd90}: color_data = 12'ha86;
			{8'd134, 8'd91}: color_data = 12'hd97;
			{8'd134, 8'd92}: color_data = 12'hc97;
			{8'd134, 8'd93}: color_data = 12'hc97;
			{8'd134, 8'd94}: color_data = 12'hc97;
			{8'd134, 8'd95}: color_data = 12'hc97;
			{8'd134, 8'd96}: color_data = 12'hc97;
			{8'd134, 8'd97}: color_data = 12'hc97;
			{8'd134, 8'd98}: color_data = 12'hc97;
			{8'd134, 8'd99}: color_data = 12'hc97;
			{8'd134, 8'd100}: color_data = 12'hc97;
			{8'd134, 8'd101}: color_data = 12'hc97;
			{8'd134, 8'd102}: color_data = 12'hc97;
			{8'd134, 8'd103}: color_data = 12'hc97;
			{8'd134, 8'd104}: color_data = 12'hc97;
			{8'd134, 8'd105}: color_data = 12'hc97;
			{8'd134, 8'd106}: color_data = 12'hc97;
			{8'd134, 8'd107}: color_data = 12'hc97;
			{8'd134, 8'd108}: color_data = 12'hc97;
			{8'd134, 8'd109}: color_data = 12'hc97;
			{8'd134, 8'd110}: color_data = 12'hc97;
			{8'd134, 8'd111}: color_data = 12'hc97;
			{8'd134, 8'd112}: color_data = 12'hc97;
			{8'd134, 8'd113}: color_data = 12'hd97;
			{8'd134, 8'd114}: color_data = 12'hc97;
			{8'd134, 8'd115}: color_data = 12'h865;
			{8'd134, 8'd116}: color_data = 12'h432;
			{8'd134, 8'd117}: color_data = 12'h000;
			{8'd135, 8'd89}: color_data = 12'h000;
			{8'd135, 8'd90}: color_data = 12'h211;
			{8'd135, 8'd91}: color_data = 12'h643;
			{8'd135, 8'd92}: color_data = 12'h975;
			{8'd135, 8'd93}: color_data = 12'hb97;
			{8'd135, 8'd94}: color_data = 12'hc97;
			{8'd135, 8'd95}: color_data = 12'hd97;
			{8'd135, 8'd96}: color_data = 12'hc97;
			{8'd135, 8'd97}: color_data = 12'hc97;
			{8'd135, 8'd98}: color_data = 12'hc97;
			{8'd135, 8'd99}: color_data = 12'hc97;
			{8'd135, 8'd100}: color_data = 12'hc97;
			{8'd135, 8'd101}: color_data = 12'hc97;
			{8'd135, 8'd102}: color_data = 12'hc97;
			{8'd135, 8'd103}: color_data = 12'hc97;
			{8'd135, 8'd104}: color_data = 12'hc97;
			{8'd135, 8'd105}: color_data = 12'hc97;
			{8'd135, 8'd106}: color_data = 12'hc97;
			{8'd135, 8'd107}: color_data = 12'hc97;
			{8'd135, 8'd108}: color_data = 12'hc97;
			{8'd135, 8'd109}: color_data = 12'hc97;
			{8'd135, 8'd110}: color_data = 12'hc97;
			{8'd135, 8'd111}: color_data = 12'hd97;
			{8'd135, 8'd112}: color_data = 12'hc97;
			{8'd135, 8'd113}: color_data = 12'h865;
			{8'd135, 8'd114}: color_data = 12'h432;
			{8'd135, 8'd115}: color_data = 12'h000;
			{8'd136, 8'd91}: color_data = 12'h000;
			{8'd136, 8'd92}: color_data = 12'h000;
			{8'd136, 8'd93}: color_data = 12'h322;
			{8'd136, 8'd94}: color_data = 12'h643;
			{8'd136, 8'd95}: color_data = 12'h864;
			{8'd136, 8'd96}: color_data = 12'h975;
			{8'd136, 8'd97}: color_data = 12'hb86;
			{8'd136, 8'd98}: color_data = 12'hc97;
			{8'd136, 8'd99}: color_data = 12'hc97;
			{8'd136, 8'd100}: color_data = 12'hd97;
			{8'd136, 8'd101}: color_data = 12'hc97;
			{8'd136, 8'd102}: color_data = 12'hc97;
			{8'd136, 8'd103}: color_data = 12'hc97;
			{8'd136, 8'd104}: color_data = 12'hc97;
			{8'd136, 8'd105}: color_data = 12'hc97;
			{8'd136, 8'd106}: color_data = 12'hc97;
			{8'd136, 8'd107}: color_data = 12'hd97;
			{8'd136, 8'd108}: color_data = 12'hd97;
			{8'd136, 8'd109}: color_data = 12'hc97;
			{8'd136, 8'd110}: color_data = 12'ha76;
			{8'd136, 8'd111}: color_data = 12'h754;
			{8'd136, 8'd112}: color_data = 12'h322;
			{8'd136, 8'd113}: color_data = 12'h000;
			{8'd137, 8'd95}: color_data = 12'h000;
			{8'd137, 8'd96}: color_data = 12'h000;
			{8'd137, 8'd97}: color_data = 12'h211;
			{8'd137, 8'd98}: color_data = 12'h432;
			{8'd137, 8'd99}: color_data = 12'h643;
			{8'd137, 8'd100}: color_data = 12'h754;
			{8'd137, 8'd101}: color_data = 12'h865;
			{8'd137, 8'd102}: color_data = 12'h976;
			{8'd137, 8'd103}: color_data = 12'hb86;
			{8'd137, 8'd104}: color_data = 12'hb87;
			{8'd137, 8'd105}: color_data = 12'ha86;
			{8'd137, 8'd106}: color_data = 12'h975;
			{8'd137, 8'd107}: color_data = 12'h865;
			{8'd137, 8'd108}: color_data = 12'h654;
			{8'd137, 8'd109}: color_data = 12'h432;
			{8'd137, 8'd110}: color_data = 12'h100;
			{8'd137, 8'd111}: color_data = 12'h000;
			{8'd138, 8'd100}: color_data = 12'h000;
			{8'd138, 8'd101}: color_data = 12'h000;
			{8'd138, 8'd102}: color_data = 12'h000;
			{8'd138, 8'd103}: color_data = 12'h211;
			{8'd138, 8'd104}: color_data = 12'h221;
			{8'd138, 8'd105}: color_data = 12'h111;
			{8'd138, 8'd106}: color_data = 12'h000;
			{8'd138, 8'd107}: color_data = 12'h000;
			{8'd138, 8'd108}: color_data = 12'h000;
            default: color_data = 12'h3b9;
        endcase
endmodule
