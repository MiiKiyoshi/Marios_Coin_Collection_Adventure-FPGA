module mario_rom_walking2(
        input wire clk,
        input wire [4:0] x,
        input wire [4:0] y,
        output reg [11:0] color_data
);

    (* rom_style = "block" *)

    //signal declaration
    reg [4:0] x_reg;
    reg [4:0] y_reg;

    always @(posedge clk) begin
        x_reg <= x;
        y_reg <= y;
    end

    always @*
        case ({x_reg, y_reg})
			// right: 5'd31, bottom: 5'd31
			{5'd0, 5'd0}: color_data = 12'h3b9;
			{5'd0, 5'd1}: color_data = 12'h3b9;
			{5'd0, 5'd2}: color_data = 12'h3b9;
			{5'd0, 5'd3}: color_data = 12'h3b9;
			{5'd0, 5'd4}: color_data = 12'h3b9;
			{5'd0, 5'd5}: color_data = 12'h3b9;
			{5'd0, 5'd6}: color_data = 12'h3b9;
			{5'd0, 5'd7}: color_data = 12'h3b9;
			{5'd0, 5'd8}: color_data = 12'h3b9;
			{5'd0, 5'd9}: color_data = 12'h3b9;
			{5'd0, 5'd10}: color_data = 12'h3b9;
			{5'd0, 5'd11}: color_data = 12'h3b9;
			{5'd0, 5'd12}: color_data = 12'h3b9;
			{5'd0, 5'd13}: color_data = 12'h3b9;
			{5'd0, 5'd14}: color_data = 12'h3b9;
			{5'd0, 5'd15}: color_data = 12'h3b9;
			{5'd0, 5'd16}: color_data = 12'hf90;
			{5'd0, 5'd17}: color_data = 12'hfa0;
			{5'd0, 5'd18}: color_data = 12'hf90;
			{5'd0, 5'd19}: color_data = 12'hf90;
			{5'd0, 5'd20}: color_data = 12'hf90;
			{5'd0, 5'd21}: color_data = 12'hf90;
			{5'd0, 5'd22}: color_data = 12'hfa1;
			{5'd0, 5'd23}: color_data = 12'h3b9;
			{5'd0, 5'd24}: color_data = 12'h3b9;
			{5'd0, 5'd25}: color_data = 12'h3b9;
			{5'd0, 5'd26}: color_data = 12'h3b9;
			{5'd0, 5'd27}: color_data = 12'h3b9;
			{5'd0, 5'd28}: color_data = 12'h3b9;
			{5'd0, 5'd29}: color_data = 12'h3b9;
			{5'd0, 5'd30}: color_data = 12'h3b9;
			{5'd0, 5'd31}: color_data = 12'h3b9;
			{5'd1, 5'd0}: color_data = 12'h3b9;
			{5'd1, 5'd1}: color_data = 12'h3b9;
			{5'd1, 5'd2}: color_data = 12'h3b9;
			{5'd1, 5'd3}: color_data = 12'h3b9;
			{5'd1, 5'd4}: color_data = 12'h3b9;
			{5'd1, 5'd5}: color_data = 12'h3b9;
			{5'd1, 5'd6}: color_data = 12'h3b9;
			{5'd1, 5'd7}: color_data = 12'h3b9;
			{5'd1, 5'd8}: color_data = 12'h3b9;
			{5'd1, 5'd9}: color_data = 12'h3b9;
			{5'd1, 5'd10}: color_data = 12'h3b9;
			{5'd1, 5'd11}: color_data = 12'h3b9;
			{5'd1, 5'd12}: color_data = 12'h3b9;
			{5'd1, 5'd13}: color_data = 12'h3b9;
			{5'd1, 5'd14}: color_data = 12'h3b9;
			{5'd1, 5'd15}: color_data = 12'h3b9;
			{5'd1, 5'd16}: color_data = 12'hfa0;
			{5'd1, 5'd17}: color_data = 12'hfa1;
			{5'd1, 5'd18}: color_data = 12'hfa1;
			{5'd1, 5'd19}: color_data = 12'hfa1;
			{5'd1, 5'd20}: color_data = 12'hfa1;
			{5'd1, 5'd21}: color_data = 12'hfa0;
			{5'd1, 5'd22}: color_data = 12'hf90;
			{5'd1, 5'd23}: color_data = 12'h3b9;
			{5'd1, 5'd24}: color_data = 12'h3b9;
			{5'd1, 5'd25}: color_data = 12'h3b9;
			{5'd1, 5'd26}: color_data = 12'h3b9;
			{5'd1, 5'd27}: color_data = 12'h3b9;
			{5'd1, 5'd28}: color_data = 12'h3b9;
			{5'd1, 5'd29}: color_data = 12'h3b9;
			{5'd1, 5'd30}: color_data = 12'h3b9;
			{5'd1, 5'd31}: color_data = 12'h3b9;
			{5'd2, 5'd0}: color_data = 12'h3b9;
			{5'd2, 5'd1}: color_data = 12'h3b9;
			{5'd2, 5'd2}: color_data = 12'h3b9;
			{5'd2, 5'd3}: color_data = 12'h3b9;
			{5'd2, 5'd4}: color_data = 12'h3b9;
			{5'd2, 5'd5}: color_data = 12'h3b9;
			{5'd2, 5'd6}: color_data = 12'h3b9;
			{5'd2, 5'd7}: color_data = 12'h3b9;
			{5'd2, 5'd8}: color_data = 12'h3b9;
			{5'd2, 5'd9}: color_data = 12'h3b9;
			{5'd2, 5'd10}: color_data = 12'h3b9;
			{5'd2, 5'd11}: color_data = 12'h3b9;
			{5'd2, 5'd12}: color_data = 12'h3b9;
			{5'd2, 5'd13}: color_data = 12'h3b9;
			{5'd2, 5'd14}: color_data = 12'h3b9;
			{5'd2, 5'd15}: color_data = 12'h3b9;
			{5'd2, 5'd16}: color_data = 12'hfa0;
			{5'd2, 5'd17}: color_data = 12'hfa1;
			{5'd2, 5'd18}: color_data = 12'hfa1;
			{5'd2, 5'd19}: color_data = 12'hfa1;
			{5'd2, 5'd20}: color_data = 12'hfa1;
			{5'd2, 5'd21}: color_data = 12'hfa0;
			{5'd2, 5'd22}: color_data = 12'hf90;
			{5'd2, 5'd23}: color_data = 12'h3b9;
			{5'd2, 5'd24}: color_data = 12'h3b9;
			{5'd2, 5'd25}: color_data = 12'h3b9;
			{5'd2, 5'd26}: color_data = 12'ha22;
			{5'd2, 5'd27}: color_data = 12'ha22;
			{5'd2, 5'd28}: color_data = 12'ha22;
			{5'd2, 5'd29}: color_data = 12'ha22;
			{5'd2, 5'd30}: color_data = 12'h933;
			{5'd2, 5'd31}: color_data = 12'h3b9;
			{5'd3, 5'd0}: color_data = 12'h3b9;
			{5'd3, 5'd1}: color_data = 12'h3b9;
			{5'd3, 5'd2}: color_data = 12'h3b9;
			{5'd3, 5'd3}: color_data = 12'h3b9;
			{5'd3, 5'd4}: color_data = 12'h3b9;
			{5'd3, 5'd5}: color_data = 12'h3b9;
			{5'd3, 5'd6}: color_data = 12'h3b9;
			{5'd3, 5'd7}: color_data = 12'h3b9;
			{5'd3, 5'd8}: color_data = 12'h3b9;
			{5'd3, 5'd9}: color_data = 12'h3b9;
			{5'd3, 5'd10}: color_data = 12'h3b9;
			{5'd3, 5'd11}: color_data = 12'h3b9;
			{5'd3, 5'd12}: color_data = 12'h3b9;
			{5'd3, 5'd13}: color_data = 12'h3b9;
			{5'd3, 5'd14}: color_data = 12'h3b9;
			{5'd3, 5'd15}: color_data = 12'h3b9;
			{5'd3, 5'd16}: color_data = 12'hfa0;
			{5'd3, 5'd17}: color_data = 12'hfa1;
			{5'd3, 5'd18}: color_data = 12'hfa1;
			{5'd3, 5'd19}: color_data = 12'hfa1;
			{5'd3, 5'd20}: color_data = 12'hfa1;
			{5'd3, 5'd21}: color_data = 12'hfa1;
			{5'd3, 5'd22}: color_data = 12'hfa0;
			{5'd3, 5'd23}: color_data = 12'h3b9;
			{5'd3, 5'd24}: color_data = 12'h3b9;
			{5'd3, 5'd25}: color_data = 12'h3b9;
			{5'd3, 5'd26}: color_data = 12'ha22;
			{5'd3, 5'd27}: color_data = 12'ha22;
			{5'd3, 5'd28}: color_data = 12'ha22;
			{5'd3, 5'd29}: color_data = 12'ha22;
			{5'd3, 5'd30}: color_data = 12'ha22;
			{5'd3, 5'd31}: color_data = 12'h3b9;
			{5'd4, 5'd0}: color_data = 12'h3b9;
			{5'd4, 5'd1}: color_data = 12'h3b9;
			{5'd4, 5'd2}: color_data = 12'h3b9;
			{5'd4, 5'd3}: color_data = 12'h3b9;
			{5'd4, 5'd4}: color_data = 12'h3b9;
			{5'd4, 5'd5}: color_data = 12'h3b9;
			{5'd4, 5'd6}: color_data = 12'h3b9;
			{5'd4, 5'd7}: color_data = 12'h3b9;
			{5'd4, 5'd8}: color_data = 12'h3b9;
			{5'd4, 5'd9}: color_data = 12'h3b9;
			{5'd4, 5'd10}: color_data = 12'h3b9;
			{5'd4, 5'd11}: color_data = 12'h3b9;
			{5'd4, 5'd12}: color_data = 12'h3b9;
			{5'd4, 5'd13}: color_data = 12'h3b9;
			{5'd4, 5'd14}: color_data = 12'ha22;
			{5'd4, 5'd15}: color_data = 12'ha22;
			{5'd4, 5'd16}: color_data = 12'hb42;
			{5'd4, 5'd17}: color_data = 12'hc52;
			{5'd4, 5'd18}: color_data = 12'hf91;
			{5'd4, 5'd19}: color_data = 12'hfa0;
			{5'd4, 5'd20}: color_data = 12'hfa0;
			{5'd4, 5'd21}: color_data = 12'hf90;
			{5'd4, 5'd22}: color_data = 12'hfb0;
			{5'd4, 5'd23}: color_data = 12'h3b9;
			{5'd4, 5'd24}: color_data = 12'hf00;
			{5'd4, 5'd25}: color_data = 12'hf00;
			{5'd4, 5'd26}: color_data = 12'ha22;
			{5'd4, 5'd27}: color_data = 12'ha22;
			{5'd4, 5'd28}: color_data = 12'ha22;
			{5'd4, 5'd29}: color_data = 12'ha22;
			{5'd4, 5'd30}: color_data = 12'ha22;
			{5'd4, 5'd31}: color_data = 12'ha22;
			{5'd5, 5'd0}: color_data = 12'h3b9;
			{5'd5, 5'd1}: color_data = 12'h3b9;
			{5'd5, 5'd2}: color_data = 12'h3b9;
			{5'd5, 5'd3}: color_data = 12'h3b9;
			{5'd5, 5'd4}: color_data = 12'h3b9;
			{5'd5, 5'd5}: color_data = 12'h3b9;
			{5'd5, 5'd6}: color_data = 12'h3b9;
			{5'd5, 5'd7}: color_data = 12'h3b9;
			{5'd5, 5'd8}: color_data = 12'h3b9;
			{5'd5, 5'd9}: color_data = 12'h3b9;
			{5'd5, 5'd10}: color_data = 12'h3b9;
			{5'd5, 5'd11}: color_data = 12'h3b9;
			{5'd5, 5'd12}: color_data = 12'h3b9;
			{5'd5, 5'd13}: color_data = 12'h3b9;
			{5'd5, 5'd14}: color_data = 12'ha22;
			{5'd5, 5'd15}: color_data = 12'ha22;
			{5'd5, 5'd16}: color_data = 12'ha22;
			{5'd5, 5'd17}: color_data = 12'ha22;
			{5'd5, 5'd18}: color_data = 12'he81;
			{5'd5, 5'd19}: color_data = 12'hfa0;
			{5'd5, 5'd20}: color_data = 12'hfa0;
			{5'd5, 5'd21}: color_data = 12'h3b9;
			{5'd5, 5'd22}: color_data = 12'h3b9;
			{5'd5, 5'd23}: color_data = 12'h3b9;
			{5'd5, 5'd24}: color_data = 12'hf00;
			{5'd5, 5'd25}: color_data = 12'hf00;
			{5'd5, 5'd26}: color_data = 12'hb22;
			{5'd5, 5'd27}: color_data = 12'h922;
			{5'd5, 5'd28}: color_data = 12'ha22;
			{5'd5, 5'd29}: color_data = 12'ha22;
			{5'd5, 5'd30}: color_data = 12'ha22;
			{5'd5, 5'd31}: color_data = 12'ha22;
			{5'd6, 5'd0}: color_data = 12'h3b9;
			{5'd6, 5'd1}: color_data = 12'h3b9;
			{5'd6, 5'd2}: color_data = 12'h3b9;
			{5'd6, 5'd3}: color_data = 12'h3b9;
			{5'd6, 5'd4}: color_data = 12'h3b9;
			{5'd6, 5'd5}: color_data = 12'h000;
			{5'd6, 5'd6}: color_data = 12'ha22;
			{5'd6, 5'd7}: color_data = 12'ha22;
			{5'd6, 5'd8}: color_data = 12'ha22;
			{5'd6, 5'd9}: color_data = 12'ha22;
			{5'd6, 5'd10}: color_data = 12'ha22;
			{5'd6, 5'd11}: color_data = 12'ha22;
			{5'd6, 5'd12}: color_data = 12'ha00;
			{5'd6, 5'd13}: color_data = 12'h3b9;
			{5'd6, 5'd14}: color_data = 12'ha22;
			{5'd6, 5'd15}: color_data = 12'ha22;
			{5'd6, 5'd16}: color_data = 12'ha22;
			{5'd6, 5'd17}: color_data = 12'ha22;
			{5'd6, 5'd18}: color_data = 12'hd71;
			{5'd6, 5'd19}: color_data = 12'hfa0;
			{5'd6, 5'd20}: color_data = 12'hf91;
			{5'd6, 5'd21}: color_data = 12'h3b9;
			{5'd6, 5'd22}: color_data = 12'hf00;
			{5'd6, 5'd23}: color_data = 12'hf00;
			{5'd6, 5'd24}: color_data = 12'hf00;
			{5'd6, 5'd25}: color_data = 12'hf00;
			{5'd6, 5'd26}: color_data = 12'he00;
			{5'd6, 5'd27}: color_data = 12'hd11;
			{5'd6, 5'd28}: color_data = 12'hb22;
			{5'd6, 5'd29}: color_data = 12'ha22;
			{5'd6, 5'd30}: color_data = 12'ha22;
			{5'd6, 5'd31}: color_data = 12'ha22;
			{5'd7, 5'd0}: color_data = 12'h3b9;
			{5'd7, 5'd1}: color_data = 12'h3b9;
			{5'd7, 5'd2}: color_data = 12'h3b9;
			{5'd7, 5'd3}: color_data = 12'h3b9;
			{5'd7, 5'd4}: color_data = 12'h3b9;
			{5'd7, 5'd5}: color_data = 12'h700;
			{5'd7, 5'd6}: color_data = 12'h912;
			{5'd7, 5'd7}: color_data = 12'ha22;
			{5'd7, 5'd8}: color_data = 12'ha22;
			{5'd7, 5'd9}: color_data = 12'ha22;
			{5'd7, 5'd10}: color_data = 12'ha22;
			{5'd7, 5'd11}: color_data = 12'ha22;
			{5'd7, 5'd12}: color_data = 12'ha11;
			{5'd7, 5'd13}: color_data = 12'h3b9;
			{5'd7, 5'd14}: color_data = 12'ha22;
			{5'd7, 5'd15}: color_data = 12'ha22;
			{5'd7, 5'd16}: color_data = 12'ha22;
			{5'd7, 5'd17}: color_data = 12'ha22;
			{5'd7, 5'd18}: color_data = 12'ha12;
			{5'd7, 5'd19}: color_data = 12'h3b9;
			{5'd7, 5'd20}: color_data = 12'h3b9;
			{5'd7, 5'd21}: color_data = 12'h3b9;
			{5'd7, 5'd22}: color_data = 12'hf00;
			{5'd7, 5'd23}: color_data = 12'hf00;
			{5'd7, 5'd24}: color_data = 12'hf00;
			{5'd7, 5'd25}: color_data = 12'hf00;
			{5'd7, 5'd26}: color_data = 12'hf00;
			{5'd7, 5'd27}: color_data = 12'hf00;
			{5'd7, 5'd28}: color_data = 12'hb11;
			{5'd7, 5'd29}: color_data = 12'ha22;
			{5'd7, 5'd30}: color_data = 12'ha22;
			{5'd7, 5'd31}: color_data = 12'ha22;
			{5'd8, 5'd0}: color_data = 12'h3b9;
			{5'd8, 5'd1}: color_data = 12'h3b9;
			{5'd8, 5'd2}: color_data = 12'hf00;
			{5'd8, 5'd3}: color_data = 12'hf00;
			{5'd8, 5'd4}: color_data = 12'ha12;
			{5'd8, 5'd5}: color_data = 12'ha22;
			{5'd8, 5'd6}: color_data = 12'hd61;
			{5'd8, 5'd7}: color_data = 12'hd61;
			{5'd8, 5'd8}: color_data = 12'hd61;
			{5'd8, 5'd9}: color_data = 12'hd61;
			{5'd8, 5'd10}: color_data = 12'ha32;
			{5'd8, 5'd11}: color_data = 12'ha22;
			{5'd8, 5'd12}: color_data = 12'ha21;
			{5'd8, 5'd13}: color_data = 12'h3b9;
			{5'd8, 5'd14}: color_data = 12'ha22;
			{5'd8, 5'd15}: color_data = 12'ha22;
			{5'd8, 5'd16}: color_data = 12'ha22;
			{5'd8, 5'd17}: color_data = 12'ha22;
			{5'd8, 5'd18}: color_data = 12'ha22;
			{5'd8, 5'd19}: color_data = 12'ha22;
			{5'd8, 5'd20}: color_data = 12'he00;
			{5'd8, 5'd21}: color_data = 12'hf00;
			{5'd8, 5'd22}: color_data = 12'hf00;
			{5'd8, 5'd23}: color_data = 12'hf00;
			{5'd8, 5'd24}: color_data = 12'hf00;
			{5'd8, 5'd25}: color_data = 12'hf00;
			{5'd8, 5'd26}: color_data = 12'hf00;
			{5'd8, 5'd27}: color_data = 12'hf00;
			{5'd8, 5'd28}: color_data = 12'hc11;
			{5'd8, 5'd29}: color_data = 12'h922;
			{5'd8, 5'd30}: color_data = 12'ha22;
			{5'd8, 5'd31}: color_data = 12'ha22;
			{5'd9, 5'd0}: color_data = 12'h3b9;
			{5'd9, 5'd1}: color_data = 12'hf00;
			{5'd9, 5'd2}: color_data = 12'hf00;
			{5'd9, 5'd3}: color_data = 12'hf00;
			{5'd9, 5'd4}: color_data = 12'hb22;
			{5'd9, 5'd5}: color_data = 12'ha22;
			{5'd9, 5'd6}: color_data = 12'hf91;
			{5'd9, 5'd7}: color_data = 12'hfa0;
			{5'd9, 5'd8}: color_data = 12'hfa0;
			{5'd9, 5'd9}: color_data = 12'hfa1;
			{5'd9, 5'd10}: color_data = 12'hb32;
			{5'd9, 5'd11}: color_data = 12'h922;
			{5'd9, 5'd12}: color_data = 12'h911;
			{5'd9, 5'd13}: color_data = 12'h3b9;
			{5'd9, 5'd14}: color_data = 12'ha22;
			{5'd9, 5'd15}: color_data = 12'ha22;
			{5'd9, 5'd16}: color_data = 12'ha22;
			{5'd9, 5'd17}: color_data = 12'ha22;
			{5'd9, 5'd18}: color_data = 12'ha22;
			{5'd9, 5'd19}: color_data = 12'ha22;
			{5'd9, 5'd20}: color_data = 12'he00;
			{5'd9, 5'd21}: color_data = 12'hf00;
			{5'd9, 5'd22}: color_data = 12'hf00;
			{5'd9, 5'd23}: color_data = 12'hf00;
			{5'd9, 5'd24}: color_data = 12'hf00;
			{5'd9, 5'd25}: color_data = 12'hf00;
			{5'd9, 5'd26}: color_data = 12'hf00;
			{5'd9, 5'd27}: color_data = 12'hf00;
			{5'd9, 5'd28}: color_data = 12'hf00;
			{5'd9, 5'd29}: color_data = 12'h3b9;
			{5'd9, 5'd30}: color_data = 12'ha22;
			{5'd9, 5'd31}: color_data = 12'ha22;
			{5'd10, 5'd0}: color_data = 12'h3b9;
			{5'd10, 5'd1}: color_data = 12'hf00;
			{5'd10, 5'd2}: color_data = 12'hf00;
			{5'd10, 5'd3}: color_data = 12'hf00;
			{5'd10, 5'd4}: color_data = 12'ha22;
			{5'd10, 5'd5}: color_data = 12'ha22;
			{5'd10, 5'd6}: color_data = 12'he81;
			{5'd10, 5'd7}: color_data = 12'hf91;
			{5'd10, 5'd8}: color_data = 12'hf91;
			{5'd10, 5'd9}: color_data = 12'hf91;
			{5'd10, 5'd10}: color_data = 12'hb42;
			{5'd10, 5'd11}: color_data = 12'ha22;
			{5'd10, 5'd12}: color_data = 12'hc41;
			{5'd10, 5'd13}: color_data = 12'h3b9;
			{5'd10, 5'd14}: color_data = 12'ha22;
			{5'd10, 5'd15}: color_data = 12'ha22;
			{5'd10, 5'd16}: color_data = 12'ha22;
			{5'd10, 5'd17}: color_data = 12'ha22;
			{5'd10, 5'd18}: color_data = 12'ha22;
			{5'd10, 5'd19}: color_data = 12'ha22;
			{5'd10, 5'd20}: color_data = 12'he00;
			{5'd10, 5'd21}: color_data = 12'hf00;
			{5'd10, 5'd22}: color_data = 12'hf00;
			{5'd10, 5'd23}: color_data = 12'hf00;
			{5'd10, 5'd24}: color_data = 12'hf00;
			{5'd10, 5'd25}: color_data = 12'hf00;
			{5'd10, 5'd26}: color_data = 12'hf00;
			{5'd10, 5'd27}: color_data = 12'hf00;
			{5'd10, 5'd28}: color_data = 12'hf00;
			{5'd10, 5'd29}: color_data = 12'h3b9;
			{5'd10, 5'd30}: color_data = 12'ha22;
			{5'd10, 5'd31}: color_data = 12'ha22;
			{5'd11, 5'd0}: color_data = 12'hf00;
			{5'd11, 5'd1}: color_data = 12'hf00;
			{5'd11, 5'd2}: color_data = 12'hf00;
			{5'd11, 5'd3}: color_data = 12'hf00;
			{5'd11, 5'd4}: color_data = 12'ha22;
			{5'd11, 5'd5}: color_data = 12'ha22;
			{5'd11, 5'd6}: color_data = 12'ha32;
			{5'd11, 5'd7}: color_data = 12'ha32;
			{5'd11, 5'd8}: color_data = 12'ha32;
			{5'd11, 5'd9}: color_data = 12'ha32;
			{5'd11, 5'd10}: color_data = 12'he81;
			{5'd11, 5'd11}: color_data = 12'hf91;
			{5'd11, 5'd12}: color_data = 12'hfa0;
			{5'd11, 5'd13}: color_data = 12'hfa0;
			{5'd11, 5'd14}: color_data = 12'ha32;
			{5'd11, 5'd15}: color_data = 12'ha22;
			{5'd11, 5'd16}: color_data = 12'ha22;
			{5'd11, 5'd17}: color_data = 12'ha22;
			{5'd11, 5'd18}: color_data = 12'ha22;
			{5'd11, 5'd19}: color_data = 12'ha22;
			{5'd11, 5'd20}: color_data = 12'he00;
			{5'd11, 5'd21}: color_data = 12'hf00;
			{5'd11, 5'd22}: color_data = 12'hf00;
			{5'd11, 5'd23}: color_data = 12'hf00;
			{5'd11, 5'd24}: color_data = 12'hf00;
			{5'd11, 5'd25}: color_data = 12'hf00;
			{5'd11, 5'd26}: color_data = 12'hf00;
			{5'd11, 5'd27}: color_data = 12'hf00;
			{5'd11, 5'd28}: color_data = 12'hf00;
			{5'd11, 5'd29}: color_data = 12'h3b9;
			{5'd11, 5'd30}: color_data = 12'h3b9;
			{5'd11, 5'd31}: color_data = 12'h3b9;
			{5'd12, 5'd0}: color_data = 12'hf00;
			{5'd12, 5'd1}: color_data = 12'hf00;
			{5'd12, 5'd2}: color_data = 12'hf00;
			{5'd12, 5'd3}: color_data = 12'hf00;
			{5'd12, 5'd4}: color_data = 12'ha22;
			{5'd12, 5'd5}: color_data = 12'ha22;
			{5'd12, 5'd6}: color_data = 12'ha22;
			{5'd12, 5'd7}: color_data = 12'ha22;
			{5'd12, 5'd8}: color_data = 12'ha22;
			{5'd12, 5'd9}: color_data = 12'ha22;
			{5'd12, 5'd10}: color_data = 12'he91;
			{5'd12, 5'd11}: color_data = 12'hfa1;
			{5'd12, 5'd12}: color_data = 12'hfa1;
			{5'd12, 5'd13}: color_data = 12'hfa1;
			{5'd12, 5'd14}: color_data = 12'hb32;
			{5'd12, 5'd15}: color_data = 12'ha22;
			{5'd12, 5'd16}: color_data = 12'ha22;
			{5'd12, 5'd17}: color_data = 12'ha22;
			{5'd12, 5'd18}: color_data = 12'ha22;
			{5'd12, 5'd19}: color_data = 12'ha22;
			{5'd12, 5'd20}: color_data = 12'he00;
			{5'd12, 5'd21}: color_data = 12'hf00;
			{5'd12, 5'd22}: color_data = 12'hf00;
			{5'd12, 5'd23}: color_data = 12'hf00;
			{5'd12, 5'd24}: color_data = 12'hf00;
			{5'd12, 5'd25}: color_data = 12'hf00;
			{5'd12, 5'd26}: color_data = 12'hf00;
			{5'd12, 5'd27}: color_data = 12'hf00;
			{5'd12, 5'd28}: color_data = 12'hf00;
			{5'd12, 5'd29}: color_data = 12'h3b9;
			{5'd12, 5'd30}: color_data = 12'h3b9;
			{5'd12, 5'd31}: color_data = 12'h3b9;
			{5'd13, 5'd0}: color_data = 12'hf00;
			{5'd13, 5'd1}: color_data = 12'hf00;
			{5'd13, 5'd2}: color_data = 12'hf00;
			{5'd13, 5'd3}: color_data = 12'hf00;
			{5'd13, 5'd4}: color_data = 12'ha22;
			{5'd13, 5'd5}: color_data = 12'ha22;
			{5'd13, 5'd6}: color_data = 12'he81;
			{5'd13, 5'd7}: color_data = 12'he91;
			{5'd13, 5'd8}: color_data = 12'ha32;
			{5'd13, 5'd9}: color_data = 12'ha22;
			{5'd13, 5'd10}: color_data = 12'he91;
			{5'd13, 5'd11}: color_data = 12'hfa1;
			{5'd13, 5'd12}: color_data = 12'hfa1;
			{5'd13, 5'd13}: color_data = 12'hfa1;
			{5'd13, 5'd14}: color_data = 12'hf20;
			{5'd13, 5'd15}: color_data = 12'hf00;
			{5'd13, 5'd16}: color_data = 12'hf00;
			{5'd13, 5'd17}: color_data = 12'hf00;
			{5'd13, 5'd18}: color_data = 12'hf00;
			{5'd13, 5'd19}: color_data = 12'hf00;
			{5'd13, 5'd20}: color_data = 12'hf00;
			{5'd13, 5'd21}: color_data = 12'hf00;
			{5'd13, 5'd22}: color_data = 12'hf00;
			{5'd13, 5'd23}: color_data = 12'hf00;
			{5'd13, 5'd24}: color_data = 12'hf00;
			{5'd13, 5'd25}: color_data = 12'hf00;
			{5'd13, 5'd26}: color_data = 12'hf00;
			{5'd13, 5'd27}: color_data = 12'hf00;
			{5'd13, 5'd28}: color_data = 12'hf00;
			{5'd13, 5'd29}: color_data = 12'h3b9;
			{5'd13, 5'd30}: color_data = 12'h3b9;
			{5'd13, 5'd31}: color_data = 12'h3b9;
			{5'd14, 5'd0}: color_data = 12'hf00;
			{5'd14, 5'd1}: color_data = 12'hf00;
			{5'd14, 5'd2}: color_data = 12'hf00;
			{5'd14, 5'd3}: color_data = 12'hf00;
			{5'd14, 5'd4}: color_data = 12'ha22;
			{5'd14, 5'd5}: color_data = 12'ha22;
			{5'd14, 5'd6}: color_data = 12'hf91;
			{5'd14, 5'd7}: color_data = 12'hfa1;
			{5'd14, 5'd8}: color_data = 12'hb32;
			{5'd14, 5'd9}: color_data = 12'ha22;
			{5'd14, 5'd10}: color_data = 12'he91;
			{5'd14, 5'd11}: color_data = 12'hfa1;
			{5'd14, 5'd12}: color_data = 12'hfa1;
			{5'd14, 5'd13}: color_data = 12'hfa1;
			{5'd14, 5'd14}: color_data = 12'hf20;
			{5'd14, 5'd15}: color_data = 12'hf00;
			{5'd14, 5'd16}: color_data = 12'hf00;
			{5'd14, 5'd17}: color_data = 12'hf00;
			{5'd14, 5'd18}: color_data = 12'hf00;
			{5'd14, 5'd19}: color_data = 12'hf00;
			{5'd14, 5'd20}: color_data = 12'hf00;
			{5'd14, 5'd21}: color_data = 12'hf00;
			{5'd14, 5'd22}: color_data = 12'hf00;
			{5'd14, 5'd23}: color_data = 12'hf00;
			{5'd14, 5'd24}: color_data = 12'hf00;
			{5'd14, 5'd25}: color_data = 12'hf00;
			{5'd14, 5'd26}: color_data = 12'hf00;
			{5'd14, 5'd27}: color_data = 12'h3b9;
			{5'd14, 5'd28}: color_data = 12'h3b9;
			{5'd14, 5'd29}: color_data = 12'h3b9;
			{5'd14, 5'd30}: color_data = 12'h3b9;
			{5'd14, 5'd31}: color_data = 12'h3b9;
			{5'd15, 5'd0}: color_data = 12'hf00;
			{5'd15, 5'd1}: color_data = 12'hf00;
			{5'd15, 5'd2}: color_data = 12'hf00;
			{5'd15, 5'd3}: color_data = 12'hf00;
			{5'd15, 5'd4}: color_data = 12'he71;
			{5'd15, 5'd5}: color_data = 12'he91;
			{5'd15, 5'd6}: color_data = 12'hfa1;
			{5'd15, 5'd7}: color_data = 12'hfa1;
			{5'd15, 5'd8}: color_data = 12'he91;
			{5'd15, 5'd9}: color_data = 12'he81;
			{5'd15, 5'd10}: color_data = 12'hfa1;
			{5'd15, 5'd11}: color_data = 12'hfa1;
			{5'd15, 5'd12}: color_data = 12'hfa1;
			{5'd15, 5'd13}: color_data = 12'hfa1;
			{5'd15, 5'd14}: color_data = 12'hf20;
			{5'd15, 5'd15}: color_data = 12'hf00;
			{5'd15, 5'd16}: color_data = 12'hf00;
			{5'd15, 5'd17}: color_data = 12'hf00;
			{5'd15, 5'd18}: color_data = 12'hf60;
			{5'd15, 5'd19}: color_data = 12'hf80;
			{5'd15, 5'd20}: color_data = 12'hf20;
			{5'd15, 5'd21}: color_data = 12'hf00;
			{5'd15, 5'd22}: color_data = 12'hf00;
			{5'd15, 5'd23}: color_data = 12'hf00;
			{5'd15, 5'd24}: color_data = 12'hf00;
			{5'd15, 5'd25}: color_data = 12'hf00;
			{5'd15, 5'd26}: color_data = 12'hf00;
			{5'd15, 5'd27}: color_data = 12'h3b9;
			{5'd15, 5'd28}: color_data = 12'h3b9;
			{5'd15, 5'd29}: color_data = 12'h3b9;
			{5'd15, 5'd30}: color_data = 12'h3b9;
			{5'd15, 5'd31}: color_data = 12'h3b9;
			{5'd16, 5'd0}: color_data = 12'hf00;
			{5'd16, 5'd1}: color_data = 12'hf00;
			{5'd16, 5'd2}: color_data = 12'hf00;
			{5'd16, 5'd3}: color_data = 12'hf00;
			{5'd16, 5'd4}: color_data = 12'hf90;
			{5'd16, 5'd5}: color_data = 12'hfa0;
			{5'd16, 5'd6}: color_data = 12'hfa1;
			{5'd16, 5'd7}: color_data = 12'hfa1;
			{5'd16, 5'd8}: color_data = 12'hfa0;
			{5'd16, 5'd9}: color_data = 12'hfa0;
			{5'd16, 5'd10}: color_data = 12'hfa1;
			{5'd16, 5'd11}: color_data = 12'hfa1;
			{5'd16, 5'd12}: color_data = 12'hfa1;
			{5'd16, 5'd13}: color_data = 12'hfa1;
			{5'd16, 5'd14}: color_data = 12'hf20;
			{5'd16, 5'd15}: color_data = 12'hf00;
			{5'd16, 5'd16}: color_data = 12'hf00;
			{5'd16, 5'd17}: color_data = 12'hf00;
			{5'd16, 5'd18}: color_data = 12'hf80;
			{5'd16, 5'd19}: color_data = 12'hfb1;
			{5'd16, 5'd20}: color_data = 12'hf20;
			{5'd16, 5'd21}: color_data = 12'hf00;
			{5'd16, 5'd22}: color_data = 12'hf00;
			{5'd16, 5'd23}: color_data = 12'hf00;
			{5'd16, 5'd24}: color_data = 12'hf00;
			{5'd16, 5'd25}: color_data = 12'hf00;
			{5'd16, 5'd26}: color_data = 12'hf00;
			{5'd16, 5'd27}: color_data = 12'h3b9;
			{5'd16, 5'd28}: color_data = 12'h3b9;
			{5'd16, 5'd29}: color_data = 12'h3b9;
			{5'd16, 5'd30}: color_data = 12'h3b9;
			{5'd16, 5'd31}: color_data = 12'h3b9;
			{5'd17, 5'd0}: color_data = 12'hf00;
			{5'd17, 5'd1}: color_data = 12'hf00;
			{5'd17, 5'd2}: color_data = 12'hf00;
			{5'd17, 5'd3}: color_data = 12'hf00;
			{5'd17, 5'd4}: color_data = 12'hf90;
			{5'd17, 5'd5}: color_data = 12'hfa1;
			{5'd17, 5'd6}: color_data = 12'hfa1;
			{5'd17, 5'd7}: color_data = 12'hfa1;
			{5'd17, 5'd8}: color_data = 12'hfa1;
			{5'd17, 5'd9}: color_data = 12'hfa1;
			{5'd17, 5'd10}: color_data = 12'hfa1;
			{5'd17, 5'd11}: color_data = 12'hfa1;
			{5'd17, 5'd12}: color_data = 12'hfa1;
			{5'd17, 5'd13}: color_data = 12'hfa1;
			{5'd17, 5'd14}: color_data = 12'hc31;
			{5'd17, 5'd15}: color_data = 12'hb12;
			{5'd17, 5'd16}: color_data = 12'hf00;
			{5'd17, 5'd17}: color_data = 12'hf00;
			{5'd17, 5'd18}: color_data = 12'hf20;
			{5'd17, 5'd19}: color_data = 12'hf20;
			{5'd17, 5'd20}: color_data = 12'hf00;
			{5'd17, 5'd21}: color_data = 12'hf00;
			{5'd17, 5'd22}: color_data = 12'hf00;
			{5'd17, 5'd23}: color_data = 12'hf00;
			{5'd17, 5'd24}: color_data = 12'hf00;
			{5'd17, 5'd25}: color_data = 12'hf00;
			{5'd17, 5'd26}: color_data = 12'hf00;
			{5'd17, 5'd27}: color_data = 12'h3b9;
			{5'd17, 5'd28}: color_data = 12'h3b9;
			{5'd17, 5'd29}: color_data = 12'h3b9;
			{5'd17, 5'd30}: color_data = 12'h3b9;
			{5'd17, 5'd31}: color_data = 12'h3b9;
			{5'd18, 5'd0}: color_data = 12'hf00;
			{5'd18, 5'd1}: color_data = 12'hf00;
			{5'd18, 5'd2}: color_data = 12'hf00;
			{5'd18, 5'd3}: color_data = 12'hf00;
			{5'd18, 5'd4}: color_data = 12'hf90;
			{5'd18, 5'd5}: color_data = 12'hfa1;
			{5'd18, 5'd6}: color_data = 12'hfa1;
			{5'd18, 5'd7}: color_data = 12'hfa1;
			{5'd18, 5'd8}: color_data = 12'hfa1;
			{5'd18, 5'd9}: color_data = 12'hfa1;
			{5'd18, 5'd10}: color_data = 12'hfa1;
			{5'd18, 5'd11}: color_data = 12'hfa1;
			{5'd18, 5'd12}: color_data = 12'hfa1;
			{5'd18, 5'd13}: color_data = 12'hfa1;
			{5'd18, 5'd14}: color_data = 12'hb42;
			{5'd18, 5'd15}: color_data = 12'h922;
			{5'd18, 5'd16}: color_data = 12'he00;
			{5'd18, 5'd17}: color_data = 12'hf00;
			{5'd18, 5'd18}: color_data = 12'hf00;
			{5'd18, 5'd19}: color_data = 12'hf00;
			{5'd18, 5'd20}: color_data = 12'hf00;
			{5'd18, 5'd21}: color_data = 12'hf00;
			{5'd18, 5'd22}: color_data = 12'hf00;
			{5'd18, 5'd23}: color_data = 12'hf00;
			{5'd18, 5'd24}: color_data = 12'hf00;
			{5'd18, 5'd25}: color_data = 12'hf00;
			{5'd18, 5'd26}: color_data = 12'hf00;
			{5'd18, 5'd27}: color_data = 12'h3b9;
			{5'd18, 5'd28}: color_data = 12'h3b9;
			{5'd18, 5'd29}: color_data = 12'h3b9;
			{5'd18, 5'd30}: color_data = 12'h3b9;
			{5'd18, 5'd31}: color_data = 12'h3b9;
			{5'd19, 5'd0}: color_data = 12'hf00;
			{5'd19, 5'd1}: color_data = 12'hf00;
			{5'd19, 5'd2}: color_data = 12'hf00;
			{5'd19, 5'd3}: color_data = 12'hf00;
			{5'd19, 5'd4}: color_data = 12'hc41;
			{5'd19, 5'd5}: color_data = 12'hb52;
			{5'd19, 5'd6}: color_data = 12'hb42;
			{5'd19, 5'd7}: color_data = 12'hc42;
			{5'd19, 5'd8}: color_data = 12'hf91;
			{5'd19, 5'd9}: color_data = 12'hfa1;
			{5'd19, 5'd10}: color_data = 12'hc51;
			{5'd19, 5'd11}: color_data = 12'hb42;
			{5'd19, 5'd12}: color_data = 12'hf91;
			{5'd19, 5'd13}: color_data = 12'hfa1;
			{5'd19, 5'd14}: color_data = 12'hb32;
			{5'd19, 5'd15}: color_data = 12'ha22;
			{5'd19, 5'd16}: color_data = 12'hb22;
			{5'd19, 5'd17}: color_data = 12'hb11;
			{5'd19, 5'd18}: color_data = 12'hf00;
			{5'd19, 5'd19}: color_data = 12'hf00;
			{5'd19, 5'd20}: color_data = 12'hf00;
			{5'd19, 5'd21}: color_data = 12'hf00;
			{5'd19, 5'd22}: color_data = 12'hf00;
			{5'd19, 5'd23}: color_data = 12'hf00;
			{5'd19, 5'd24}: color_data = 12'hf00;
			{5'd19, 5'd25}: color_data = 12'hf00;
			{5'd19, 5'd26}: color_data = 12'hf00;
			{5'd19, 5'd27}: color_data = 12'hf00;
			{5'd19, 5'd28}: color_data = 12'hf00;
			{5'd19, 5'd29}: color_data = 12'h3b9;
			{5'd19, 5'd30}: color_data = 12'h3b9;
			{5'd19, 5'd31}: color_data = 12'h3b9;
			{5'd20, 5'd0}: color_data = 12'hf00;
			{5'd20, 5'd1}: color_data = 12'hf00;
			{5'd20, 5'd2}: color_data = 12'hf00;
			{5'd20, 5'd3}: color_data = 12'hf00;
			{5'd20, 5'd4}: color_data = 12'ha12;
			{5'd20, 5'd5}: color_data = 12'h922;
			{5'd20, 5'd6}: color_data = 12'h912;
			{5'd20, 5'd7}: color_data = 12'h922;
			{5'd20, 5'd8}: color_data = 12'hf91;
			{5'd20, 5'd9}: color_data = 12'hfa0;
			{5'd20, 5'd10}: color_data = 12'ha32;
			{5'd20, 5'd11}: color_data = 12'ha22;
			{5'd20, 5'd12}: color_data = 12'he91;
			{5'd20, 5'd13}: color_data = 12'hfa1;
			{5'd20, 5'd14}: color_data = 12'hb32;
			{5'd20, 5'd15}: color_data = 12'ha22;
			{5'd20, 5'd16}: color_data = 12'ha22;
			{5'd20, 5'd17}: color_data = 12'ha22;
			{5'd20, 5'd18}: color_data = 12'he00;
			{5'd20, 5'd19}: color_data = 12'hf00;
			{5'd20, 5'd20}: color_data = 12'hf00;
			{5'd20, 5'd21}: color_data = 12'hf00;
			{5'd20, 5'd22}: color_data = 12'hf00;
			{5'd20, 5'd23}: color_data = 12'hf00;
			{5'd20, 5'd24}: color_data = 12'hf00;
			{5'd20, 5'd25}: color_data = 12'hf00;
			{5'd20, 5'd26}: color_data = 12'hf00;
			{5'd20, 5'd27}: color_data = 12'hf00;
			{5'd20, 5'd28}: color_data = 12'hf00;
			{5'd20, 5'd29}: color_data = 12'h3b9;
			{5'd20, 5'd30}: color_data = 12'h3b9;
			{5'd20, 5'd31}: color_data = 12'h3b9;
			{5'd21, 5'd0}: color_data = 12'hf00;
			{5'd21, 5'd1}: color_data = 12'hf00;
			{5'd21, 5'd2}: color_data = 12'hf00;
			{5'd21, 5'd3}: color_data = 12'hf00;
			{5'd21, 5'd4}: color_data = 12'he61;
			{5'd21, 5'd5}: color_data = 12'hd71;
			{5'd21, 5'd6}: color_data = 12'hd71;
			{5'd21, 5'd7}: color_data = 12'hd71;
			{5'd21, 5'd8}: color_data = 12'hc51;
			{5'd21, 5'd9}: color_data = 12'hc52;
			{5'd21, 5'd10}: color_data = 12'ha22;
			{5'd21, 5'd11}: color_data = 12'ha22;
			{5'd21, 5'd12}: color_data = 12'he91;
			{5'd21, 5'd13}: color_data = 12'hfa0;
			{5'd21, 5'd14}: color_data = 12'hd61;
			{5'd21, 5'd15}: color_data = 12'h902;
			{5'd21, 5'd16}: color_data = 12'ha22;
			{5'd21, 5'd17}: color_data = 12'ha22;
			{5'd21, 5'd18}: color_data = 12'he00;
			{5'd21, 5'd19}: color_data = 12'hf00;
			{5'd21, 5'd20}: color_data = 12'hf00;
			{5'd21, 5'd21}: color_data = 12'hf00;
			{5'd21, 5'd22}: color_data = 12'hf00;
			{5'd21, 5'd23}: color_data = 12'hf00;
			{5'd21, 5'd24}: color_data = 12'hf00;
			{5'd21, 5'd25}: color_data = 12'hf00;
			{5'd21, 5'd26}: color_data = 12'hf00;
			{5'd21, 5'd27}: color_data = 12'hf00;
			{5'd21, 5'd28}: color_data = 12'hf00;
			{5'd21, 5'd29}: color_data = 12'h3b9;
			{5'd21, 5'd30}: color_data = 12'h3b9;
			{5'd21, 5'd31}: color_data = 12'h3b9;
			{5'd22, 5'd0}: color_data = 12'h3b9;
			{5'd22, 5'd1}: color_data = 12'h3b9;
			{5'd22, 5'd2}: color_data = 12'hf00;
			{5'd22, 5'd3}: color_data = 12'hf00;
			{5'd22, 5'd4}: color_data = 12'hf90;
			{5'd22, 5'd5}: color_data = 12'hfa0;
			{5'd22, 5'd6}: color_data = 12'hfa0;
			{5'd22, 5'd7}: color_data = 12'hfa1;
			{5'd22, 5'd8}: color_data = 12'ha32;
			{5'd22, 5'd9}: color_data = 12'h912;
			{5'd22, 5'd10}: color_data = 12'ha22;
			{5'd22, 5'd11}: color_data = 12'ha22;
			{5'd22, 5'd12}: color_data = 12'hf91;
			{5'd22, 5'd13}: color_data = 12'hfa0;
			{5'd22, 5'd14}: color_data = 12'hf90;
			{5'd22, 5'd15}: color_data = 12'h3b9;
			{5'd22, 5'd16}: color_data = 12'ha22;
			{5'd22, 5'd17}: color_data = 12'ha22;
			{5'd22, 5'd18}: color_data = 12'he00;
			{5'd22, 5'd19}: color_data = 12'hf00;
			{5'd22, 5'd20}: color_data = 12'hf00;
			{5'd22, 5'd21}: color_data = 12'hf00;
			{5'd22, 5'd22}: color_data = 12'hf00;
			{5'd22, 5'd23}: color_data = 12'hf00;
			{5'd22, 5'd24}: color_data = 12'hf00;
			{5'd22, 5'd25}: color_data = 12'hf00;
			{5'd22, 5'd26}: color_data = 12'hf00;
			{5'd22, 5'd27}: color_data = 12'hf00;
			{5'd22, 5'd28}: color_data = 12'hf00;
			{5'd22, 5'd29}: color_data = 12'h3b9;
			{5'd22, 5'd30}: color_data = 12'h3b9;
			{5'd22, 5'd31}: color_data = 12'h3b9;
			{5'd23, 5'd0}: color_data = 12'h3b9;
			{5'd23, 5'd1}: color_data = 12'hf00;
			{5'd23, 5'd2}: color_data = 12'hf00;
			{5'd23, 5'd3}: color_data = 12'hf00;
			{5'd23, 5'd4}: color_data = 12'hf70;
			{5'd23, 5'd5}: color_data = 12'hfa0;
			{5'd23, 5'd6}: color_data = 12'hfa0;
			{5'd23, 5'd7}: color_data = 12'hfa1;
			{5'd23, 5'd8}: color_data = 12'hd71;
			{5'd23, 5'd9}: color_data = 12'hd61;
			{5'd23, 5'd10}: color_data = 12'ha32;
			{5'd23, 5'd11}: color_data = 12'ha22;
			{5'd23, 5'd12}: color_data = 12'hf91;
			{5'd23, 5'd13}: color_data = 12'hfa0;
			{5'd23, 5'd14}: color_data = 12'hf90;
			{5'd23, 5'd15}: color_data = 12'h3b9;
			{5'd23, 5'd16}: color_data = 12'ha22;
			{5'd23, 5'd17}: color_data = 12'ha22;
			{5'd23, 5'd18}: color_data = 12'hc11;
			{5'd23, 5'd19}: color_data = 12'hc11;
			{5'd23, 5'd20}: color_data = 12'he00;
			{5'd23, 5'd21}: color_data = 12'hf00;
			{5'd23, 5'd22}: color_data = 12'hf00;
			{5'd23, 5'd23}: color_data = 12'hf00;
			{5'd23, 5'd24}: color_data = 12'hf00;
			{5'd23, 5'd25}: color_data = 12'hf00;
			{5'd23, 5'd26}: color_data = 12'hf00;
			{5'd23, 5'd27}: color_data = 12'hf00;
			{5'd23, 5'd28}: color_data = 12'hf00;
			{5'd23, 5'd29}: color_data = 12'h3b9;
			{5'd23, 5'd30}: color_data = 12'h3b9;
			{5'd23, 5'd31}: color_data = 12'h3b9;
			{5'd24, 5'd0}: color_data = 12'h3b9;
			{5'd24, 5'd1}: color_data = 12'hf00;
			{5'd24, 5'd2}: color_data = 12'hf00;
			{5'd24, 5'd3}: color_data = 12'hf00;
			{5'd24, 5'd4}: color_data = 12'hf00;
			{5'd24, 5'd5}: color_data = 12'h3b9;
			{5'd24, 5'd6}: color_data = 12'hfa0;
			{5'd24, 5'd7}: color_data = 12'hfa1;
			{5'd24, 5'd8}: color_data = 12'hfa0;
			{5'd24, 5'd9}: color_data = 12'hfa1;
			{5'd24, 5'd10}: color_data = 12'hb32;
			{5'd24, 5'd11}: color_data = 12'ha22;
			{5'd24, 5'd12}: color_data = 12'hf91;
			{5'd24, 5'd13}: color_data = 12'hfa0;
			{5'd24, 5'd14}: color_data = 12'hf90;
			{5'd24, 5'd15}: color_data = 12'h3b9;
			{5'd24, 5'd16}: color_data = 12'h922;
			{5'd24, 5'd17}: color_data = 12'ha22;
			{5'd24, 5'd18}: color_data = 12'ha22;
			{5'd24, 5'd19}: color_data = 12'h922;
			{5'd24, 5'd20}: color_data = 12'h922;
			{5'd24, 5'd21}: color_data = 12'h3b9;
			{5'd24, 5'd22}: color_data = 12'hf00;
			{5'd24, 5'd23}: color_data = 12'hf00;
			{5'd24, 5'd24}: color_data = 12'hf00;
			{5'd24, 5'd25}: color_data = 12'hf00;
			{5'd24, 5'd26}: color_data = 12'hf00;
			{5'd24, 5'd27}: color_data = 12'hf00;
			{5'd24, 5'd28}: color_data = 12'hf00;
			{5'd24, 5'd29}: color_data = 12'h3b9;
			{5'd24, 5'd30}: color_data = 12'h3b9;
			{5'd24, 5'd31}: color_data = 12'h3b9;
			{5'd25, 5'd0}: color_data = 12'h3b9;
			{5'd25, 5'd1}: color_data = 12'hf00;
			{5'd25, 5'd2}: color_data = 12'hf00;
			{5'd25, 5'd3}: color_data = 12'hf00;
			{5'd25, 5'd4}: color_data = 12'hf00;
			{5'd25, 5'd5}: color_data = 12'h3b9;
			{5'd25, 5'd6}: color_data = 12'hfa0;
			{5'd25, 5'd7}: color_data = 12'hfa1;
			{5'd25, 5'd8}: color_data = 12'hfa1;
			{5'd25, 5'd9}: color_data = 12'hfa1;
			{5'd25, 5'd10}: color_data = 12'hb32;
			{5'd25, 5'd11}: color_data = 12'ha22;
			{5'd25, 5'd12}: color_data = 12'he71;
			{5'd25, 5'd13}: color_data = 12'hfa0;
			{5'd25, 5'd14}: color_data = 12'hfa1;
			{5'd25, 5'd15}: color_data = 12'h3b9;
			{5'd25, 5'd16}: color_data = 12'hd61;
			{5'd25, 5'd17}: color_data = 12'hd61;
			{5'd25, 5'd18}: color_data = 12'ha32;
			{5'd25, 5'd19}: color_data = 12'ha22;
			{5'd25, 5'd20}: color_data = 12'h921;
			{5'd25, 5'd21}: color_data = 12'h3b9;
			{5'd25, 5'd22}: color_data = 12'hc11;
			{5'd25, 5'd23}: color_data = 12'hd11;
			{5'd25, 5'd24}: color_data = 12'hc11;
			{5'd25, 5'd25}: color_data = 12'hc11;
			{5'd25, 5'd26}: color_data = 12'hd11;
			{5'd25, 5'd27}: color_data = 12'hc11;
			{5'd25, 5'd28}: color_data = 12'hc00;
			{5'd25, 5'd29}: color_data = 12'h3b9;
			{5'd25, 5'd30}: color_data = 12'h3b9;
			{5'd25, 5'd31}: color_data = 12'h3b9;
			{5'd26, 5'd0}: color_data = 12'h3b9;
			{5'd26, 5'd1}: color_data = 12'hf00;
			{5'd26, 5'd2}: color_data = 12'hf00;
			{5'd26, 5'd3}: color_data = 12'hf00;
			{5'd26, 5'd4}: color_data = 12'hf00;
			{5'd26, 5'd5}: color_data = 12'hff0;
			{5'd26, 5'd6}: color_data = 12'hfa0;
			{5'd26, 5'd7}: color_data = 12'hfa1;
			{5'd26, 5'd8}: color_data = 12'hfa1;
			{5'd26, 5'd9}: color_data = 12'hfa1;
			{5'd26, 5'd10}: color_data = 12'hb32;
			{5'd26, 5'd11}: color_data = 12'ha22;
			{5'd26, 5'd12}: color_data = 12'h911;
			{5'd26, 5'd13}: color_data = 12'h3b9;
			{5'd26, 5'd14}: color_data = 12'h3b9;
			{5'd26, 5'd15}: color_data = 12'h3b9;
			{5'd26, 5'd16}: color_data = 12'hfa0;
			{5'd26, 5'd17}: color_data = 12'hfb1;
			{5'd26, 5'd18}: color_data = 12'hb32;
			{5'd26, 5'd19}: color_data = 12'h912;
			{5'd26, 5'd20}: color_data = 12'h911;
			{5'd26, 5'd21}: color_data = 12'h3b9;
			{5'd26, 5'd22}: color_data = 12'h922;
			{5'd26, 5'd23}: color_data = 12'ha22;
			{5'd26, 5'd24}: color_data = 12'ha22;
			{5'd26, 5'd25}: color_data = 12'ha22;
			{5'd26, 5'd26}: color_data = 12'ha22;
			{5'd26, 5'd27}: color_data = 12'h922;
			{5'd26, 5'd28}: color_data = 12'h911;
			{5'd26, 5'd29}: color_data = 12'h3b9;
			{5'd26, 5'd30}: color_data = 12'h3b9;
			{5'd26, 5'd31}: color_data = 12'h3b9;
			{5'd27, 5'd0}: color_data = 12'h3b9;
			{5'd27, 5'd1}: color_data = 12'h3b9;
			{5'd27, 5'd2}: color_data = 12'hf00;
			{5'd27, 5'd3}: color_data = 12'hf00;
			{5'd27, 5'd4}: color_data = 12'hf00;
			{5'd27, 5'd5}: color_data = 12'h3b9;
			{5'd27, 5'd6}: color_data = 12'hf91;
			{5'd27, 5'd7}: color_data = 12'hf90;
			{5'd27, 5'd8}: color_data = 12'hfa1;
			{5'd27, 5'd9}: color_data = 12'hfa0;
			{5'd27, 5'd10}: color_data = 12'hb41;
			{5'd27, 5'd11}: color_data = 12'h912;
			{5'd27, 5'd12}: color_data = 12'ha00;
			{5'd27, 5'd13}: color_data = 12'h3b9;
			{5'd27, 5'd14}: color_data = 12'h3b9;
			{5'd27, 5'd15}: color_data = 12'h3b9;
			{5'd27, 5'd16}: color_data = 12'hfa0;
			{5'd27, 5'd17}: color_data = 12'hfa1;
			{5'd27, 5'd18}: color_data = 12'hd61;
			{5'd27, 5'd19}: color_data = 12'hc51;
			{5'd27, 5'd20}: color_data = 12'hb41;
			{5'd27, 5'd21}: color_data = 12'ha12;
			{5'd27, 5'd22}: color_data = 12'ha22;
			{5'd27, 5'd23}: color_data = 12'ha22;
			{5'd27, 5'd24}: color_data = 12'ha22;
			{5'd27, 5'd25}: color_data = 12'ha22;
			{5'd27, 5'd26}: color_data = 12'ha22;
			{5'd27, 5'd27}: color_data = 12'ha22;
			{5'd27, 5'd28}: color_data = 12'ha11;
			{5'd27, 5'd29}: color_data = 12'h3b9;
			{5'd27, 5'd30}: color_data = 12'h3b9;
			{5'd27, 5'd31}: color_data = 12'h3b9;
			{5'd28, 5'd0}: color_data = 12'h3b9;
			{5'd28, 5'd1}: color_data = 12'h3b9;
			{5'd28, 5'd2}: color_data = 12'h3b9;
			{5'd28, 5'd3}: color_data = 12'h3b9;
			{5'd28, 5'd4}: color_data = 12'h3b9;
			{5'd28, 5'd5}: color_data = 12'h3b9;
			{5'd28, 5'd6}: color_data = 12'h3b9;
			{5'd28, 5'd7}: color_data = 12'hfa0;
			{5'd28, 5'd8}: color_data = 12'hfa0;
			{5'd28, 5'd9}: color_data = 12'hfa1;
			{5'd28, 5'd10}: color_data = 12'hfa1;
			{5'd28, 5'd11}: color_data = 12'h3b9;
			{5'd28, 5'd12}: color_data = 12'h3b9;
			{5'd28, 5'd13}: color_data = 12'h3b9;
			{5'd28, 5'd14}: color_data = 12'h3b9;
			{5'd28, 5'd15}: color_data = 12'h3b9;
			{5'd28, 5'd16}: color_data = 12'hfa0;
			{5'd28, 5'd17}: color_data = 12'hfa1;
			{5'd28, 5'd18}: color_data = 12'hfa0;
			{5'd28, 5'd19}: color_data = 12'hfa0;
			{5'd28, 5'd20}: color_data = 12'hb42;
			{5'd28, 5'd21}: color_data = 12'ha22;
			{5'd28, 5'd22}: color_data = 12'ha22;
			{5'd28, 5'd23}: color_data = 12'ha22;
			{5'd28, 5'd24}: color_data = 12'ha22;
			{5'd28, 5'd25}: color_data = 12'ha22;
			{5'd28, 5'd26}: color_data = 12'ha22;
			{5'd28, 5'd27}: color_data = 12'ha22;
			{5'd28, 5'd28}: color_data = 12'ha11;
			{5'd28, 5'd29}: color_data = 12'h3b9;
			{5'd28, 5'd30}: color_data = 12'h3b9;
			{5'd28, 5'd31}: color_data = 12'h3b9;
			{5'd29, 5'd0}: color_data = 12'h3b9;
			{5'd29, 5'd1}: color_data = 12'h3b9;
			{5'd29, 5'd2}: color_data = 12'h3b9;
			{5'd29, 5'd3}: color_data = 12'h3b9;
			{5'd29, 5'd4}: color_data = 12'h3b9;
			{5'd29, 5'd5}: color_data = 12'h3b9;
			{5'd29, 5'd6}: color_data = 12'h3b9;
			{5'd29, 5'd7}: color_data = 12'hff0;
			{5'd29, 5'd8}: color_data = 12'hf90;
			{5'd29, 5'd9}: color_data = 12'hf90;
			{5'd29, 5'd10}: color_data = 12'hf70;
			{5'd29, 5'd11}: color_data = 12'h3b9;
			{5'd29, 5'd12}: color_data = 12'h3b9;
			{5'd29, 5'd13}: color_data = 12'h3b9;
			{5'd29, 5'd14}: color_data = 12'h3b9;
			{5'd29, 5'd15}: color_data = 12'h3b9;
			{5'd29, 5'd16}: color_data = 12'hfa0;
			{5'd29, 5'd17}: color_data = 12'hfa1;
			{5'd29, 5'd18}: color_data = 12'hfa1;
			{5'd29, 5'd19}: color_data = 12'hfa0;
			{5'd29, 5'd20}: color_data = 12'hc51;
			{5'd29, 5'd21}: color_data = 12'h912;
			{5'd29, 5'd22}: color_data = 12'ha22;
			{5'd29, 5'd23}: color_data = 12'ha22;
			{5'd29, 5'd24}: color_data = 12'ha22;
			{5'd29, 5'd25}: color_data = 12'ha22;
			{5'd29, 5'd26}: color_data = 12'ha22;
			{5'd29, 5'd27}: color_data = 12'h922;
			{5'd29, 5'd28}: color_data = 12'ha22;
			{5'd29, 5'd29}: color_data = 12'h3b9;
			{5'd29, 5'd30}: color_data = 12'h3b9;
			{5'd29, 5'd31}: color_data = 12'h3b9;
			{5'd30, 5'd0}: color_data = 12'h3b9;
			{5'd30, 5'd1}: color_data = 12'h3b9;
			{5'd30, 5'd2}: color_data = 12'h3b9;
			{5'd30, 5'd3}: color_data = 12'h3b9;
			{5'd30, 5'd4}: color_data = 12'h3b9;
			{5'd30, 5'd5}: color_data = 12'h3b9;
			{5'd30, 5'd6}: color_data = 12'h3b9;
			{5'd30, 5'd7}: color_data = 12'h3b9;
			{5'd30, 5'd8}: color_data = 12'h3b9;
			{5'd30, 5'd9}: color_data = 12'h3b9;
			{5'd30, 5'd10}: color_data = 12'h3b9;
			{5'd30, 5'd11}: color_data = 12'h3b9;
			{5'd30, 5'd12}: color_data = 12'h3b9;
			{5'd30, 5'd13}: color_data = 12'h3b9;
			{5'd30, 5'd14}: color_data = 12'h3b9;
			{5'd30, 5'd15}: color_data = 12'h3b9;
			{5'd30, 5'd16}: color_data = 12'hfa0;
			{5'd30, 5'd17}: color_data = 12'hfa1;
			{5'd30, 5'd18}: color_data = 12'hfa1;
			{5'd30, 5'd19}: color_data = 12'hfa0;
			{5'd30, 5'd20}: color_data = 12'hfa0;
			{5'd30, 5'd21}: color_data = 12'h3b9;
			{5'd30, 5'd22}: color_data = 12'h3b9;
			{5'd30, 5'd23}: color_data = 12'h3b9;
			{5'd30, 5'd24}: color_data = 12'h3b9;
			{5'd30, 5'd25}: color_data = 12'h3b9;
			{5'd30, 5'd26}: color_data = 12'h3b9;
			{5'd30, 5'd27}: color_data = 12'h3b9;
			{5'd30, 5'd28}: color_data = 12'h3b9;
			{5'd30, 5'd29}: color_data = 12'h3b9;
			{5'd30, 5'd30}: color_data = 12'h3b9;
			{5'd30, 5'd31}: color_data = 12'h3b9;
			{5'd31, 5'd0}: color_data = 12'h3b9;
			{5'd31, 5'd1}: color_data = 12'h3b9;
			{5'd31, 5'd2}: color_data = 12'h3b9;
			{5'd31, 5'd3}: color_data = 12'h3b9;
			{5'd31, 5'd4}: color_data = 12'h3b9;
			{5'd31, 5'd5}: color_data = 12'h3b9;
			{5'd31, 5'd6}: color_data = 12'h3b9;
			{5'd31, 5'd7}: color_data = 12'h3b9;
			{5'd31, 5'd8}: color_data = 12'h3b9;
			{5'd31, 5'd9}: color_data = 12'h3b9;
			{5'd31, 5'd10}: color_data = 12'h3b9;
			{5'd31, 5'd11}: color_data = 12'h3b9;
			{5'd31, 5'd12}: color_data = 12'h3b9;
			{5'd31, 5'd13}: color_data = 12'h3b9;
			{5'd31, 5'd14}: color_data = 12'h3b9;
			{5'd31, 5'd15}: color_data = 12'h3b9;
			{5'd31, 5'd16}: color_data = 12'hf90;
			{5'd31, 5'd17}: color_data = 12'hf90;
			{5'd31, 5'd18}: color_data = 12'hf90;
			{5'd31, 5'd19}: color_data = 12'hf90;
			{5'd31, 5'd20}: color_data = 12'hf91;
			{5'd31, 5'd21}: color_data = 12'h3b9;
			{5'd31, 5'd22}: color_data = 12'h3b9;
			{5'd31, 5'd23}: color_data = 12'h3b9;
			{5'd31, 5'd24}: color_data = 12'h3b9;
			{5'd31, 5'd25}: color_data = 12'h3b9;
			{5'd31, 5'd26}: color_data = 12'h3b9;
			{5'd31, 5'd27}: color_data = 12'h3b9;
			{5'd31, 5'd28}: color_data = 12'h3b9;
			{5'd31, 5'd29}: color_data = 12'h3b9;
			{5'd31, 5'd30}: color_data = 12'h3b9;
			{5'd31, 5'd31}: color_data = 12'h3b9;
            default: color_data = 12'h3b9;
        endcase
endmodule
