module goomba_rom(
        input wire clk,
        input wire [4:0] x,
        input wire [4:0] y,
        output reg [11:0] color_data
);

    (* rom_style = "block" *)

    //signal declaration
    reg [4:0] x_reg;
    reg [4:0] y_reg;

    always @(posedge clk) begin
        x_reg <= x;
        y_reg <= y;
    end

    always @*
        case ({x_reg, y_reg})
			// right: 5'd26, bottom: 5'd27
			{5'd0, 5'd0}: color_data = 12'h3b9;
			{5'd0, 5'd1}: color_data = 12'h3b9;
			{5'd0, 5'd2}: color_data = 12'h3b9;
			{5'd0, 5'd3}: color_data = 12'h3b9;
			{5'd0, 5'd4}: color_data = 12'h3b9;
			{5'd0, 5'd5}: color_data = 12'h3b9;
			{5'd0, 5'd6}: color_data = 12'h3b9;
			{5'd0, 5'd7}: color_data = 12'h3b9;
			{5'd0, 5'd8}: color_data = 12'h3b9;
			{5'd0, 5'd9}: color_data = 12'h3b9;
			{5'd0, 5'd10}: color_data = 12'h3b9;
			{5'd0, 5'd11}: color_data = 12'h3b9;
			{5'd0, 5'd12}: color_data = 12'h752;
			{5'd0, 5'd13}: color_data = 12'h752;
			{5'd0, 5'd14}: color_data = 12'h742;
			{5'd0, 5'd15}: color_data = 12'h742;
			{5'd0, 5'd16}: color_data = 12'h752;
			{5'd0, 5'd17}: color_data = 12'h752;
			{5'd0, 5'd18}: color_data = 12'h3b9;
			{5'd0, 5'd19}: color_data = 12'h3b9;
			{5'd0, 5'd20}: color_data = 12'h3b9;
			{5'd0, 5'd21}: color_data = 12'h3b9;
			{5'd0, 5'd22}: color_data = 12'h3b9;
			{5'd0, 5'd23}: color_data = 12'h3b9;
			{5'd0, 5'd24}: color_data = 12'h3b9;
			{5'd0, 5'd25}: color_data = 12'h3b9;
			{5'd0, 5'd26}: color_data = 12'h3b9;
			{5'd0, 5'd27}: color_data = 12'h3b9;
			{5'd1, 5'd0}: color_data = 12'h3b9;
			{5'd1, 5'd1}: color_data = 12'h3b9;
			{5'd1, 5'd2}: color_data = 12'h3b9;
			{5'd1, 5'd3}: color_data = 12'h3b9;
			{5'd1, 5'd4}: color_data = 12'h3b9;
			{5'd1, 5'd5}: color_data = 12'h3b9;
			{5'd1, 5'd6}: color_data = 12'h3b9;
			{5'd1, 5'd7}: color_data = 12'h3b9;
			{5'd1, 5'd8}: color_data = 12'h853;
			{5'd1, 5'd9}: color_data = 12'h752;
			{5'd1, 5'd10}: color_data = 12'h752;
			{5'd1, 5'd11}: color_data = 12'h752;
			{5'd1, 5'd12}: color_data = 12'h752;
			{5'd1, 5'd13}: color_data = 12'h752;
			{5'd1, 5'd14}: color_data = 12'h752;
			{5'd1, 5'd15}: color_data = 12'h752;
			{5'd1, 5'd16}: color_data = 12'h752;
			{5'd1, 5'd17}: color_data = 12'h752;
			{5'd1, 5'd18}: color_data = 12'h752;
			{5'd1, 5'd19}: color_data = 12'h852;
			{5'd1, 5'd20}: color_data = 12'h3b9;
			{5'd1, 5'd21}: color_data = 12'h3b9;
			{5'd1, 5'd22}: color_data = 12'h000;
			{5'd1, 5'd23}: color_data = 12'h000;
			{5'd1, 5'd24}: color_data = 12'h000;
			{5'd1, 5'd25}: color_data = 12'h000;
			{5'd1, 5'd26}: color_data = 12'h000;
			{5'd1, 5'd27}: color_data = 12'h3b9;
			{5'd2, 5'd0}: color_data = 12'h3b9;
			{5'd2, 5'd1}: color_data = 12'h3b9;
			{5'd2, 5'd2}: color_data = 12'h3b9;
			{5'd2, 5'd3}: color_data = 12'h3b9;
			{5'd2, 5'd4}: color_data = 12'h3b9;
			{5'd2, 5'd5}: color_data = 12'h3b9;
			{5'd2, 5'd6}: color_data = 12'h3b9;
			{5'd2, 5'd7}: color_data = 12'h3b9;
			{5'd2, 5'd8}: color_data = 12'h752;
			{5'd2, 5'd9}: color_data = 12'h752;
			{5'd2, 5'd10}: color_data = 12'h752;
			{5'd2, 5'd11}: color_data = 12'h752;
			{5'd2, 5'd12}: color_data = 12'h752;
			{5'd2, 5'd13}: color_data = 12'h752;
			{5'd2, 5'd14}: color_data = 12'h752;
			{5'd2, 5'd15}: color_data = 12'h752;
			{5'd2, 5'd16}: color_data = 12'h752;
			{5'd2, 5'd17}: color_data = 12'h752;
			{5'd2, 5'd18}: color_data = 12'h852;
			{5'd2, 5'd19}: color_data = 12'h752;
			{5'd2, 5'd20}: color_data = 12'h3b9;
			{5'd2, 5'd21}: color_data = 12'h3b9;
			{5'd2, 5'd22}: color_data = 12'h000;
			{5'd2, 5'd23}: color_data = 12'h000;
			{5'd2, 5'd24}: color_data = 12'h000;
			{5'd2, 5'd25}: color_data = 12'h000;
			{5'd2, 5'd26}: color_data = 12'h000;
			{5'd2, 5'd27}: color_data = 12'h3b9;
			{5'd3, 5'd0}: color_data = 12'h3b9;
			{5'd3, 5'd1}: color_data = 12'h3b9;
			{5'd3, 5'd2}: color_data = 12'h3b9;
			{5'd3, 5'd3}: color_data = 12'h3b9;
			{5'd3, 5'd4}: color_data = 12'h3b9;
			{5'd3, 5'd5}: color_data = 12'h3b9;
			{5'd3, 5'd6}: color_data = 12'h752;
			{5'd3, 5'd7}: color_data = 12'h752;
			{5'd3, 5'd8}: color_data = 12'h752;
			{5'd3, 5'd9}: color_data = 12'h742;
			{5'd3, 5'd10}: color_data = 12'h752;
			{5'd3, 5'd11}: color_data = 12'h752;
			{5'd3, 5'd12}: color_data = 12'h752;
			{5'd3, 5'd13}: color_data = 12'h752;
			{5'd3, 5'd14}: color_data = 12'h752;
			{5'd3, 5'd15}: color_data = 12'h752;
			{5'd3, 5'd16}: color_data = 12'h752;
			{5'd3, 5'd17}: color_data = 12'h752;
			{5'd3, 5'd18}: color_data = 12'h752;
			{5'd3, 5'd19}: color_data = 12'h752;
			{5'd3, 5'd20}: color_data = 12'h000;
			{5'd3, 5'd21}: color_data = 12'h000;
			{5'd3, 5'd22}: color_data = 12'h000;
			{5'd3, 5'd23}: color_data = 12'h000;
			{5'd3, 5'd24}: color_data = 12'h000;
			{5'd3, 5'd25}: color_data = 12'h000;
			{5'd3, 5'd26}: color_data = 12'h000;
			{5'd3, 5'd27}: color_data = 12'h000;
			{5'd4, 5'd0}: color_data = 12'h3b9;
			{5'd4, 5'd1}: color_data = 12'h3b9;
			{5'd4, 5'd2}: color_data = 12'h3b9;
			{5'd4, 5'd3}: color_data = 12'h3b9;
			{5'd4, 5'd4}: color_data = 12'h3b9;
			{5'd4, 5'd5}: color_data = 12'h752;
			{5'd4, 5'd6}: color_data = 12'h752;
			{5'd4, 5'd7}: color_data = 12'h742;
			{5'd4, 5'd8}: color_data = 12'h752;
			{5'd4, 5'd9}: color_data = 12'h752;
			{5'd4, 5'd10}: color_data = 12'h752;
			{5'd4, 5'd11}: color_data = 12'h752;
			{5'd4, 5'd12}: color_data = 12'h752;
			{5'd4, 5'd13}: color_data = 12'h752;
			{5'd4, 5'd14}: color_data = 12'h752;
			{5'd4, 5'd15}: color_data = 12'h752;
			{5'd4, 5'd16}: color_data = 12'h752;
			{5'd4, 5'd17}: color_data = 12'h752;
			{5'd4, 5'd18}: color_data = 12'h752;
			{5'd4, 5'd19}: color_data = 12'h852;
			{5'd4, 5'd20}: color_data = 12'h000;
			{5'd4, 5'd21}: color_data = 12'h000;
			{5'd4, 5'd22}: color_data = 12'h000;
			{5'd4, 5'd23}: color_data = 12'h000;
			{5'd4, 5'd24}: color_data = 12'h000;
			{5'd4, 5'd25}: color_data = 12'h000;
			{5'd4, 5'd26}: color_data = 12'h000;
			{5'd4, 5'd27}: color_data = 12'h000;
			{5'd5, 5'd0}: color_data = 12'h3b9;
			{5'd5, 5'd1}: color_data = 12'h3b9;
			{5'd5, 5'd2}: color_data = 12'h3b9;
			{5'd5, 5'd3}: color_data = 12'h3b9;
			{5'd5, 5'd4}: color_data = 12'h3b9;
			{5'd5, 5'd5}: color_data = 12'h752;
			{5'd5, 5'd6}: color_data = 12'h742;
			{5'd5, 5'd7}: color_data = 12'h100;
			{5'd5, 5'd8}: color_data = 12'h210;
			{5'd5, 5'd9}: color_data = 12'h742;
			{5'd5, 5'd10}: color_data = 12'h742;
			{5'd5, 5'd11}: color_data = 12'h742;
			{5'd5, 5'd12}: color_data = 12'h742;
			{5'd5, 5'd13}: color_data = 12'h742;
			{5'd5, 5'd14}: color_data = 12'h742;
			{5'd5, 5'd15}: color_data = 12'h742;
			{5'd5, 5'd16}: color_data = 12'h752;
			{5'd5, 5'd17}: color_data = 12'h752;
			{5'd5, 5'd18}: color_data = 12'h752;
			{5'd5, 5'd19}: color_data = 12'h752;
			{5'd5, 5'd20}: color_data = 12'h000;
			{5'd5, 5'd21}: color_data = 12'h000;
			{5'd5, 5'd22}: color_data = 12'h000;
			{5'd5, 5'd23}: color_data = 12'h000;
			{5'd5, 5'd24}: color_data = 12'h000;
			{5'd5, 5'd25}: color_data = 12'h000;
			{5'd5, 5'd26}: color_data = 12'h000;
			{5'd5, 5'd27}: color_data = 12'h000;
			{5'd6, 5'd0}: color_data = 12'h3b9;
			{5'd6, 5'd1}: color_data = 12'h3b9;
			{5'd6, 5'd2}: color_data = 12'h3b9;
			{5'd6, 5'd3}: color_data = 12'h752;
			{5'd6, 5'd4}: color_data = 12'h752;
			{5'd6, 5'd5}: color_data = 12'h752;
			{5'd6, 5'd6}: color_data = 12'h752;
			{5'd6, 5'd7}: color_data = 12'h000;
			{5'd6, 5'd8}: color_data = 12'h111;
			{5'd6, 5'd9}: color_data = 12'h986;
			{5'd6, 5'd10}: color_data = 12'h986;
			{5'd6, 5'd11}: color_data = 12'h986;
			{5'd6, 5'd12}: color_data = 12'h986;
			{5'd6, 5'd13}: color_data = 12'h986;
			{5'd6, 5'd14}: color_data = 12'h986;
			{5'd6, 5'd15}: color_data = 12'h975;
			{5'd6, 5'd16}: color_data = 12'h742;
			{5'd6, 5'd17}: color_data = 12'h752;
			{5'd6, 5'd18}: color_data = 12'h752;
			{5'd6, 5'd19}: color_data = 12'hb95;
			{5'd6, 5'd20}: color_data = 12'hdb7;
			{5'd6, 5'd21}: color_data = 12'h542;
			{5'd6, 5'd22}: color_data = 12'h321;
			{5'd6, 5'd23}: color_data = 12'h000;
			{5'd6, 5'd24}: color_data = 12'h000;
			{5'd6, 5'd25}: color_data = 12'h000;
			{5'd6, 5'd26}: color_data = 12'h000;
			{5'd6, 5'd27}: color_data = 12'h000;
			{5'd7, 5'd0}: color_data = 12'h3b9;
			{5'd7, 5'd1}: color_data = 12'h3b9;
			{5'd7, 5'd2}: color_data = 12'h3b9;
			{5'd7, 5'd3}: color_data = 12'h752;
			{5'd7, 5'd4}: color_data = 12'h752;
			{5'd7, 5'd5}: color_data = 12'h752;
			{5'd7, 5'd6}: color_data = 12'h742;
			{5'd7, 5'd7}: color_data = 12'h000;
			{5'd7, 5'd8}: color_data = 12'h333;
			{5'd7, 5'd9}: color_data = 12'hfff;
			{5'd7, 5'd10}: color_data = 12'hfff;
			{5'd7, 5'd11}: color_data = 12'hfff;
			{5'd7, 5'd12}: color_data = 12'hfff;
			{5'd7, 5'd13}: color_data = 12'hfff;
			{5'd7, 5'd14}: color_data = 12'hfff;
			{5'd7, 5'd15}: color_data = 12'hddc;
			{5'd7, 5'd16}: color_data = 12'h742;
			{5'd7, 5'd17}: color_data = 12'h742;
			{5'd7, 5'd18}: color_data = 12'h642;
			{5'd7, 5'd19}: color_data = 12'hda6;
			{5'd7, 5'd20}: color_data = 12'hfd8;
			{5'd7, 5'd21}: color_data = 12'hfd8;
			{5'd7, 5'd22}: color_data = 12'hb96;
			{5'd7, 5'd23}: color_data = 12'h000;
			{5'd7, 5'd24}: color_data = 12'h000;
			{5'd7, 5'd25}: color_data = 12'h000;
			{5'd7, 5'd26}: color_data = 12'h000;
			{5'd7, 5'd27}: color_data = 12'h000;
			{5'd8, 5'd0}: color_data = 12'h3b9;
			{5'd8, 5'd1}: color_data = 12'h742;
			{5'd8, 5'd2}: color_data = 12'h742;
			{5'd8, 5'd3}: color_data = 12'h742;
			{5'd8, 5'd4}: color_data = 12'h752;
			{5'd8, 5'd5}: color_data = 12'h752;
			{5'd8, 5'd6}: color_data = 12'h742;
			{5'd8, 5'd7}: color_data = 12'h431;
			{5'd8, 5'd8}: color_data = 12'h432;
			{5'd8, 5'd9}: color_data = 12'h666;
			{5'd8, 5'd10}: color_data = 12'h666;
			{5'd8, 5'd11}: color_data = 12'h666;
			{5'd8, 5'd12}: color_data = 12'h666;
			{5'd8, 5'd13}: color_data = 12'h777;
			{5'd8, 5'd14}: color_data = 12'hfff;
			{5'd8, 5'd15}: color_data = 12'hedc;
			{5'd8, 5'd16}: color_data = 12'h742;
			{5'd8, 5'd17}: color_data = 12'h974;
			{5'd8, 5'd18}: color_data = 12'hc95;
			{5'd8, 5'd19}: color_data = 12'heb7;
			{5'd8, 5'd20}: color_data = 12'hfc8;
			{5'd8, 5'd21}: color_data = 12'hfc8;
			{5'd8, 5'd22}: color_data = 12'hb96;
			{5'd8, 5'd23}: color_data = 12'h000;
			{5'd8, 5'd24}: color_data = 12'h000;
			{5'd8, 5'd25}: color_data = 12'h000;
			{5'd8, 5'd26}: color_data = 12'h000;
			{5'd8, 5'd27}: color_data = 12'h000;
			{5'd9, 5'd0}: color_data = 12'h3b9;
			{5'd9, 5'd1}: color_data = 12'h742;
			{5'd9, 5'd2}: color_data = 12'h752;
			{5'd9, 5'd3}: color_data = 12'h752;
			{5'd9, 5'd4}: color_data = 12'h752;
			{5'd9, 5'd5}: color_data = 12'h752;
			{5'd9, 5'd6}: color_data = 12'h752;
			{5'd9, 5'd7}: color_data = 12'h752;
			{5'd9, 5'd8}: color_data = 12'h642;
			{5'd9, 5'd9}: color_data = 12'h000;
			{5'd9, 5'd10}: color_data = 12'h000;
			{5'd9, 5'd11}: color_data = 12'h000;
			{5'd9, 5'd12}: color_data = 12'h000;
			{5'd9, 5'd13}: color_data = 12'h000;
			{5'd9, 5'd14}: color_data = 12'heee;
			{5'd9, 5'd15}: color_data = 12'hedc;
			{5'd9, 5'd16}: color_data = 12'h742;
			{5'd9, 5'd17}: color_data = 12'hb85;
			{5'd9, 5'd18}: color_data = 12'hfd8;
			{5'd9, 5'd19}: color_data = 12'hfc8;
			{5'd9, 5'd20}: color_data = 12'hfc8;
			{5'd9, 5'd21}: color_data = 12'hfc8;
			{5'd9, 5'd22}: color_data = 12'hb96;
			{5'd9, 5'd23}: color_data = 12'h000;
			{5'd9, 5'd24}: color_data = 12'h000;
			{5'd9, 5'd25}: color_data = 12'h000;
			{5'd9, 5'd26}: color_data = 12'h000;
			{5'd9, 5'd27}: color_data = 12'h000;
			{5'd10, 5'd0}: color_data = 12'h752;
			{5'd10, 5'd1}: color_data = 12'h742;
			{5'd10, 5'd2}: color_data = 12'h752;
			{5'd10, 5'd3}: color_data = 12'h752;
			{5'd10, 5'd4}: color_data = 12'h752;
			{5'd10, 5'd5}: color_data = 12'h752;
			{5'd10, 5'd6}: color_data = 12'h752;
			{5'd10, 5'd7}: color_data = 12'h752;
			{5'd10, 5'd8}: color_data = 12'h742;
			{5'd10, 5'd9}: color_data = 12'h642;
			{5'd10, 5'd10}: color_data = 12'h321;
			{5'd10, 5'd11}: color_data = 12'h000;
			{5'd10, 5'd12}: color_data = 12'h999;
			{5'd10, 5'd13}: color_data = 12'heee;
			{5'd10, 5'd14}: color_data = 12'hfff;
			{5'd10, 5'd15}: color_data = 12'hddc;
			{5'd10, 5'd16}: color_data = 12'h742;
			{5'd10, 5'd17}: color_data = 12'hb85;
			{5'd10, 5'd18}: color_data = 12'hfc8;
			{5'd10, 5'd19}: color_data = 12'hfc8;
			{5'd10, 5'd20}: color_data = 12'hfc8;
			{5'd10, 5'd21}: color_data = 12'hfc8;
			{5'd10, 5'd22}: color_data = 12'hfc7;
			{5'd10, 5'd23}: color_data = 12'hdb7;
			{5'd10, 5'd24}: color_data = 12'h653;
			{5'd10, 5'd25}: color_data = 12'h000;
			{5'd10, 5'd26}: color_data = 12'h000;
			{5'd10, 5'd27}: color_data = 12'h000;
			{5'd11, 5'd0}: color_data = 12'h752;
			{5'd11, 5'd1}: color_data = 12'h752;
			{5'd11, 5'd2}: color_data = 12'h752;
			{5'd11, 5'd3}: color_data = 12'h752;
			{5'd11, 5'd4}: color_data = 12'h752;
			{5'd11, 5'd5}: color_data = 12'h752;
			{5'd11, 5'd6}: color_data = 12'h752;
			{5'd11, 5'd7}: color_data = 12'h752;
			{5'd11, 5'd8}: color_data = 12'h752;
			{5'd11, 5'd9}: color_data = 12'h752;
			{5'd11, 5'd10}: color_data = 12'h421;
			{5'd11, 5'd11}: color_data = 12'h000;
			{5'd11, 5'd12}: color_data = 12'h999;
			{5'd11, 5'd13}: color_data = 12'heed;
			{5'd11, 5'd14}: color_data = 12'hedd;
			{5'd11, 5'd15}: color_data = 12'hcba;
			{5'd11, 5'd16}: color_data = 12'h742;
			{5'd11, 5'd17}: color_data = 12'hb85;
			{5'd11, 5'd18}: color_data = 12'hfc8;
			{5'd11, 5'd19}: color_data = 12'hfc8;
			{5'd11, 5'd20}: color_data = 12'hfc8;
			{5'd11, 5'd21}: color_data = 12'hfc8;
			{5'd11, 5'd22}: color_data = 12'hfc8;
			{5'd11, 5'd23}: color_data = 12'hfd8;
			{5'd11, 5'd24}: color_data = 12'h975;
			{5'd11, 5'd25}: color_data = 12'h321;
			{5'd11, 5'd26}: color_data = 12'h110;
			{5'd11, 5'd27}: color_data = 12'h000;
			{5'd12, 5'd0}: color_data = 12'h752;
			{5'd12, 5'd1}: color_data = 12'h752;
			{5'd12, 5'd2}: color_data = 12'h752;
			{5'd12, 5'd3}: color_data = 12'h752;
			{5'd12, 5'd4}: color_data = 12'h752;
			{5'd12, 5'd5}: color_data = 12'h752;
			{5'd12, 5'd6}: color_data = 12'h752;
			{5'd12, 5'd7}: color_data = 12'h752;
			{5'd12, 5'd8}: color_data = 12'h752;
			{5'd12, 5'd9}: color_data = 12'h752;
			{5'd12, 5'd10}: color_data = 12'h421;
			{5'd12, 5'd11}: color_data = 12'h000;
			{5'd12, 5'd12}: color_data = 12'h531;
			{5'd12, 5'd13}: color_data = 12'h752;
			{5'd12, 5'd14}: color_data = 12'h742;
			{5'd12, 5'd15}: color_data = 12'h742;
			{5'd12, 5'd16}: color_data = 12'h742;
			{5'd12, 5'd17}: color_data = 12'hb85;
			{5'd12, 5'd18}: color_data = 12'hfc8;
			{5'd12, 5'd19}: color_data = 12'hfc8;
			{5'd12, 5'd20}: color_data = 12'hfc8;
			{5'd12, 5'd21}: color_data = 12'hfc8;
			{5'd12, 5'd22}: color_data = 12'hfc8;
			{5'd12, 5'd23}: color_data = 12'hfc8;
			{5'd12, 5'd24}: color_data = 12'hfc8;
			{5'd12, 5'd25}: color_data = 12'hfc8;
			{5'd12, 5'd26}: color_data = 12'heb7;
			{5'd12, 5'd27}: color_data = 12'h000;
			{5'd13, 5'd0}: color_data = 12'h752;
			{5'd13, 5'd1}: color_data = 12'h752;
			{5'd13, 5'd2}: color_data = 12'h752;
			{5'd13, 5'd3}: color_data = 12'h752;
			{5'd13, 5'd4}: color_data = 12'h752;
			{5'd13, 5'd5}: color_data = 12'h752;
			{5'd13, 5'd6}: color_data = 12'h752;
			{5'd13, 5'd7}: color_data = 12'h752;
			{5'd13, 5'd8}: color_data = 12'h752;
			{5'd13, 5'd9}: color_data = 12'h752;
			{5'd13, 5'd10}: color_data = 12'h421;
			{5'd13, 5'd11}: color_data = 12'h000;
			{5'd13, 5'd12}: color_data = 12'h531;
			{5'd13, 5'd13}: color_data = 12'h752;
			{5'd13, 5'd14}: color_data = 12'h742;
			{5'd13, 5'd15}: color_data = 12'h742;
			{5'd13, 5'd16}: color_data = 12'h742;
			{5'd13, 5'd17}: color_data = 12'hb85;
			{5'd13, 5'd18}: color_data = 12'hfc8;
			{5'd13, 5'd19}: color_data = 12'hfc8;
			{5'd13, 5'd20}: color_data = 12'hfc8;
			{5'd13, 5'd21}: color_data = 12'hfc8;
			{5'd13, 5'd22}: color_data = 12'hfc8;
			{5'd13, 5'd23}: color_data = 12'hfc8;
			{5'd13, 5'd24}: color_data = 12'hfc8;
			{5'd13, 5'd25}: color_data = 12'hfc8;
			{5'd13, 5'd26}: color_data = 12'hfc8;
			{5'd13, 5'd27}: color_data = 12'h3b9;
			{5'd14, 5'd0}: color_data = 12'h752;
			{5'd14, 5'd1}: color_data = 12'h752;
			{5'd14, 5'd2}: color_data = 12'h752;
			{5'd14, 5'd3}: color_data = 12'h752;
			{5'd14, 5'd4}: color_data = 12'h752;
			{5'd14, 5'd5}: color_data = 12'h752;
			{5'd14, 5'd6}: color_data = 12'h752;
			{5'd14, 5'd7}: color_data = 12'h752;
			{5'd14, 5'd8}: color_data = 12'h752;
			{5'd14, 5'd9}: color_data = 12'h752;
			{5'd14, 5'd10}: color_data = 12'h421;
			{5'd14, 5'd11}: color_data = 12'h000;
			{5'd14, 5'd12}: color_data = 12'h531;
			{5'd14, 5'd13}: color_data = 12'h752;
			{5'd14, 5'd14}: color_data = 12'h742;
			{5'd14, 5'd15}: color_data = 12'h742;
			{5'd14, 5'd16}: color_data = 12'h742;
			{5'd14, 5'd17}: color_data = 12'hb85;
			{5'd14, 5'd18}: color_data = 12'hfc8;
			{5'd14, 5'd19}: color_data = 12'hfc8;
			{5'd14, 5'd20}: color_data = 12'hfc8;
			{5'd14, 5'd21}: color_data = 12'hfc8;
			{5'd14, 5'd22}: color_data = 12'hfc8;
			{5'd14, 5'd23}: color_data = 12'hfc8;
			{5'd14, 5'd24}: color_data = 12'hfc8;
			{5'd14, 5'd25}: color_data = 12'hfc8;
			{5'd14, 5'd26}: color_data = 12'heb7;
			{5'd14, 5'd27}: color_data = 12'h000;
			{5'd15, 5'd0}: color_data = 12'h752;
			{5'd15, 5'd1}: color_data = 12'h752;
			{5'd15, 5'd2}: color_data = 12'h752;
			{5'd15, 5'd3}: color_data = 12'h752;
			{5'd15, 5'd4}: color_data = 12'h752;
			{5'd15, 5'd5}: color_data = 12'h752;
			{5'd15, 5'd6}: color_data = 12'h752;
			{5'd15, 5'd7}: color_data = 12'h752;
			{5'd15, 5'd8}: color_data = 12'h752;
			{5'd15, 5'd9}: color_data = 12'h752;
			{5'd15, 5'd10}: color_data = 12'h421;
			{5'd15, 5'd11}: color_data = 12'h000;
			{5'd15, 5'd12}: color_data = 12'h999;
			{5'd15, 5'd13}: color_data = 12'heed;
			{5'd15, 5'd14}: color_data = 12'hedd;
			{5'd15, 5'd15}: color_data = 12'hcba;
			{5'd15, 5'd16}: color_data = 12'h742;
			{5'd15, 5'd17}: color_data = 12'hb85;
			{5'd15, 5'd18}: color_data = 12'hfc8;
			{5'd15, 5'd19}: color_data = 12'hfc8;
			{5'd15, 5'd20}: color_data = 12'hfc8;
			{5'd15, 5'd21}: color_data = 12'hfc8;
			{5'd15, 5'd22}: color_data = 12'hfc8;
			{5'd15, 5'd23}: color_data = 12'hfd8;
			{5'd15, 5'd24}: color_data = 12'h975;
			{5'd15, 5'd25}: color_data = 12'h221;
			{5'd15, 5'd26}: color_data = 12'h110;
			{5'd15, 5'd27}: color_data = 12'h000;
			{5'd16, 5'd0}: color_data = 12'h752;
			{5'd16, 5'd1}: color_data = 12'h752;
			{5'd16, 5'd2}: color_data = 12'h742;
			{5'd16, 5'd3}: color_data = 12'h752;
			{5'd16, 5'd4}: color_data = 12'h752;
			{5'd16, 5'd5}: color_data = 12'h752;
			{5'd16, 5'd6}: color_data = 12'h752;
			{5'd16, 5'd7}: color_data = 12'h752;
			{5'd16, 5'd8}: color_data = 12'h742;
			{5'd16, 5'd9}: color_data = 12'h642;
			{5'd16, 5'd10}: color_data = 12'h321;
			{5'd16, 5'd11}: color_data = 12'h000;
			{5'd16, 5'd12}: color_data = 12'h999;
			{5'd16, 5'd13}: color_data = 12'heee;
			{5'd16, 5'd14}: color_data = 12'hfff;
			{5'd16, 5'd15}: color_data = 12'hddc;
			{5'd16, 5'd16}: color_data = 12'h742;
			{5'd16, 5'd17}: color_data = 12'hb85;
			{5'd16, 5'd18}: color_data = 12'hfc8;
			{5'd16, 5'd19}: color_data = 12'hfc8;
			{5'd16, 5'd20}: color_data = 12'hfc8;
			{5'd16, 5'd21}: color_data = 12'hfc8;
			{5'd16, 5'd22}: color_data = 12'hfc7;
			{5'd16, 5'd23}: color_data = 12'hdb7;
			{5'd16, 5'd24}: color_data = 12'h653;
			{5'd16, 5'd25}: color_data = 12'h000;
			{5'd16, 5'd26}: color_data = 12'h000;
			{5'd16, 5'd27}: color_data = 12'h000;
			{5'd17, 5'd0}: color_data = 12'h3b9;
			{5'd17, 5'd1}: color_data = 12'h752;
			{5'd17, 5'd2}: color_data = 12'h752;
			{5'd17, 5'd3}: color_data = 12'h752;
			{5'd17, 5'd4}: color_data = 12'h752;
			{5'd17, 5'd5}: color_data = 12'h752;
			{5'd17, 5'd6}: color_data = 12'h752;
			{5'd17, 5'd7}: color_data = 12'h752;
			{5'd17, 5'd8}: color_data = 12'h642;
			{5'd17, 5'd9}: color_data = 12'h000;
			{5'd17, 5'd10}: color_data = 12'h000;
			{5'd17, 5'd11}: color_data = 12'h000;
			{5'd17, 5'd12}: color_data = 12'h000;
			{5'd17, 5'd13}: color_data = 12'h000;
			{5'd17, 5'd14}: color_data = 12'heee;
			{5'd17, 5'd15}: color_data = 12'hedc;
			{5'd17, 5'd16}: color_data = 12'h742;
			{5'd17, 5'd17}: color_data = 12'hb85;
			{5'd17, 5'd18}: color_data = 12'hfd8;
			{5'd17, 5'd19}: color_data = 12'hfc8;
			{5'd17, 5'd20}: color_data = 12'hfc8;
			{5'd17, 5'd21}: color_data = 12'hfc8;
			{5'd17, 5'd22}: color_data = 12'hb96;
			{5'd17, 5'd23}: color_data = 12'h000;
			{5'd17, 5'd24}: color_data = 12'h000;
			{5'd17, 5'd25}: color_data = 12'h000;
			{5'd17, 5'd26}: color_data = 12'h000;
			{5'd17, 5'd27}: color_data = 12'h000;
			{5'd18, 5'd0}: color_data = 12'h3b9;
			{5'd18, 5'd1}: color_data = 12'h752;
			{5'd18, 5'd2}: color_data = 12'h752;
			{5'd18, 5'd3}: color_data = 12'h752;
			{5'd18, 5'd4}: color_data = 12'h752;
			{5'd18, 5'd5}: color_data = 12'h752;
			{5'd18, 5'd6}: color_data = 12'h742;
			{5'd18, 5'd7}: color_data = 12'h431;
			{5'd18, 5'd8}: color_data = 12'h432;
			{5'd18, 5'd9}: color_data = 12'h666;
			{5'd18, 5'd10}: color_data = 12'h666;
			{5'd18, 5'd11}: color_data = 12'h666;
			{5'd18, 5'd12}: color_data = 12'h666;
			{5'd18, 5'd13}: color_data = 12'h777;
			{5'd18, 5'd14}: color_data = 12'hfff;
			{5'd18, 5'd15}: color_data = 12'hedc;
			{5'd18, 5'd16}: color_data = 12'h742;
			{5'd18, 5'd17}: color_data = 12'h974;
			{5'd18, 5'd18}: color_data = 12'hc95;
			{5'd18, 5'd19}: color_data = 12'heb7;
			{5'd18, 5'd20}: color_data = 12'hfc8;
			{5'd18, 5'd21}: color_data = 12'hfc8;
			{5'd18, 5'd22}: color_data = 12'hb96;
			{5'd18, 5'd23}: color_data = 12'h000;
			{5'd18, 5'd24}: color_data = 12'h000;
			{5'd18, 5'd25}: color_data = 12'h000;
			{5'd18, 5'd26}: color_data = 12'h000;
			{5'd18, 5'd27}: color_data = 12'h000;
			{5'd19, 5'd0}: color_data = 12'h3b9;
			{5'd19, 5'd1}: color_data = 12'h3b9;
			{5'd19, 5'd2}: color_data = 12'h3b9;
			{5'd19, 5'd3}: color_data = 12'h752;
			{5'd19, 5'd4}: color_data = 12'h752;
			{5'd19, 5'd5}: color_data = 12'h752;
			{5'd19, 5'd6}: color_data = 12'h742;
			{5'd19, 5'd7}: color_data = 12'h000;
			{5'd19, 5'd8}: color_data = 12'h333;
			{5'd19, 5'd9}: color_data = 12'hfff;
			{5'd19, 5'd10}: color_data = 12'hfff;
			{5'd19, 5'd11}: color_data = 12'hfff;
			{5'd19, 5'd12}: color_data = 12'hfff;
			{5'd19, 5'd13}: color_data = 12'hfff;
			{5'd19, 5'd14}: color_data = 12'hfff;
			{5'd19, 5'd15}: color_data = 12'hddc;
			{5'd19, 5'd16}: color_data = 12'h742;
			{5'd19, 5'd17}: color_data = 12'h742;
			{5'd19, 5'd18}: color_data = 12'h642;
			{5'd19, 5'd19}: color_data = 12'hda6;
			{5'd19, 5'd20}: color_data = 12'hfd8;
			{5'd19, 5'd21}: color_data = 12'hfd8;
			{5'd19, 5'd22}: color_data = 12'hb96;
			{5'd19, 5'd23}: color_data = 12'h000;
			{5'd19, 5'd24}: color_data = 12'h000;
			{5'd19, 5'd25}: color_data = 12'h000;
			{5'd19, 5'd26}: color_data = 12'h000;
			{5'd19, 5'd27}: color_data = 12'h000;
			{5'd20, 5'd0}: color_data = 12'h3b9;
			{5'd20, 5'd1}: color_data = 12'h3b9;
			{5'd20, 5'd2}: color_data = 12'h3b9;
			{5'd20, 5'd3}: color_data = 12'h742;
			{5'd20, 5'd4}: color_data = 12'h752;
			{5'd20, 5'd5}: color_data = 12'h752;
			{5'd20, 5'd6}: color_data = 12'h752;
			{5'd20, 5'd7}: color_data = 12'h000;
			{5'd20, 5'd8}: color_data = 12'h111;
			{5'd20, 5'd9}: color_data = 12'h976;
			{5'd20, 5'd10}: color_data = 12'h976;
			{5'd20, 5'd11}: color_data = 12'h976;
			{5'd20, 5'd12}: color_data = 12'h976;
			{5'd20, 5'd13}: color_data = 12'h976;
			{5'd20, 5'd14}: color_data = 12'h976;
			{5'd20, 5'd15}: color_data = 12'h975;
			{5'd20, 5'd16}: color_data = 12'h742;
			{5'd20, 5'd17}: color_data = 12'h752;
			{5'd20, 5'd18}: color_data = 12'h752;
			{5'd20, 5'd19}: color_data = 12'hb95;
			{5'd20, 5'd20}: color_data = 12'hdb7;
			{5'd20, 5'd21}: color_data = 12'h542;
			{5'd20, 5'd22}: color_data = 12'h321;
			{5'd20, 5'd23}: color_data = 12'h000;
			{5'd20, 5'd24}: color_data = 12'h000;
			{5'd20, 5'd25}: color_data = 12'h000;
			{5'd20, 5'd26}: color_data = 12'h000;
			{5'd20, 5'd27}: color_data = 12'h000;
			{5'd21, 5'd0}: color_data = 12'h3b9;
			{5'd21, 5'd1}: color_data = 12'h3b9;
			{5'd21, 5'd2}: color_data = 12'h3b9;
			{5'd21, 5'd3}: color_data = 12'h3b9;
			{5'd21, 5'd4}: color_data = 12'h3b9;
			{5'd21, 5'd5}: color_data = 12'h752;
			{5'd21, 5'd6}: color_data = 12'h742;
			{5'd21, 5'd7}: color_data = 12'h110;
			{5'd21, 5'd8}: color_data = 12'h210;
			{5'd21, 5'd9}: color_data = 12'h742;
			{5'd21, 5'd10}: color_data = 12'h742;
			{5'd21, 5'd11}: color_data = 12'h742;
			{5'd21, 5'd12}: color_data = 12'h742;
			{5'd21, 5'd13}: color_data = 12'h742;
			{5'd21, 5'd14}: color_data = 12'h742;
			{5'd21, 5'd15}: color_data = 12'h742;
			{5'd21, 5'd16}: color_data = 12'h752;
			{5'd21, 5'd17}: color_data = 12'h752;
			{5'd21, 5'd18}: color_data = 12'h752;
			{5'd21, 5'd19}: color_data = 12'h752;
			{5'd21, 5'd20}: color_data = 12'h000;
			{5'd21, 5'd21}: color_data = 12'h000;
			{5'd21, 5'd22}: color_data = 12'h000;
			{5'd21, 5'd23}: color_data = 12'h000;
			{5'd21, 5'd24}: color_data = 12'h000;
			{5'd21, 5'd25}: color_data = 12'h000;
			{5'd21, 5'd26}: color_data = 12'h000;
			{5'd21, 5'd27}: color_data = 12'h000;
			{5'd22, 5'd0}: color_data = 12'h3b9;
			{5'd22, 5'd1}: color_data = 12'h3b9;
			{5'd22, 5'd2}: color_data = 12'h3b9;
			{5'd22, 5'd3}: color_data = 12'h3b9;
			{5'd22, 5'd4}: color_data = 12'h3b9;
			{5'd22, 5'd5}: color_data = 12'h733;
			{5'd22, 5'd6}: color_data = 12'h752;
			{5'd22, 5'd7}: color_data = 12'h742;
			{5'd22, 5'd8}: color_data = 12'h752;
			{5'd22, 5'd9}: color_data = 12'h752;
			{5'd22, 5'd10}: color_data = 12'h752;
			{5'd22, 5'd11}: color_data = 12'h752;
			{5'd22, 5'd12}: color_data = 12'h752;
			{5'd22, 5'd13}: color_data = 12'h752;
			{5'd22, 5'd14}: color_data = 12'h752;
			{5'd22, 5'd15}: color_data = 12'h752;
			{5'd22, 5'd16}: color_data = 12'h752;
			{5'd22, 5'd17}: color_data = 12'h752;
			{5'd22, 5'd18}: color_data = 12'h752;
			{5'd22, 5'd19}: color_data = 12'h852;
			{5'd22, 5'd20}: color_data = 12'h000;
			{5'd22, 5'd21}: color_data = 12'h000;
			{5'd22, 5'd22}: color_data = 12'h000;
			{5'd22, 5'd23}: color_data = 12'h000;
			{5'd22, 5'd24}: color_data = 12'h000;
			{5'd22, 5'd25}: color_data = 12'h000;
			{5'd22, 5'd26}: color_data = 12'h000;
			{5'd22, 5'd27}: color_data = 12'h000;
			{5'd23, 5'd0}: color_data = 12'h3b9;
			{5'd23, 5'd1}: color_data = 12'h3b9;
			{5'd23, 5'd2}: color_data = 12'h3b9;
			{5'd23, 5'd3}: color_data = 12'h3b9;
			{5'd23, 5'd4}: color_data = 12'h3b9;
			{5'd23, 5'd5}: color_data = 12'h3b9;
			{5'd23, 5'd6}: color_data = 12'h752;
			{5'd23, 5'd7}: color_data = 12'h752;
			{5'd23, 5'd8}: color_data = 12'h752;
			{5'd23, 5'd9}: color_data = 12'h752;
			{5'd23, 5'd10}: color_data = 12'h752;
			{5'd23, 5'd11}: color_data = 12'h752;
			{5'd23, 5'd12}: color_data = 12'h752;
			{5'd23, 5'd13}: color_data = 12'h752;
			{5'd23, 5'd14}: color_data = 12'h752;
			{5'd23, 5'd15}: color_data = 12'h752;
			{5'd23, 5'd16}: color_data = 12'h752;
			{5'd23, 5'd17}: color_data = 12'h752;
			{5'd23, 5'd18}: color_data = 12'h752;
			{5'd23, 5'd19}: color_data = 12'h752;
			{5'd23, 5'd20}: color_data = 12'h000;
			{5'd23, 5'd21}: color_data = 12'h000;
			{5'd23, 5'd22}: color_data = 12'h000;
			{5'd23, 5'd23}: color_data = 12'h000;
			{5'd23, 5'd24}: color_data = 12'h000;
			{5'd23, 5'd25}: color_data = 12'h000;
			{5'd23, 5'd26}: color_data = 12'h000;
			{5'd23, 5'd27}: color_data = 12'h000;
			{5'd24, 5'd0}: color_data = 12'h3b9;
			{5'd24, 5'd1}: color_data = 12'h3b9;
			{5'd24, 5'd2}: color_data = 12'h3b9;
			{5'd24, 5'd3}: color_data = 12'h3b9;
			{5'd24, 5'd4}: color_data = 12'h3b9;
			{5'd24, 5'd5}: color_data = 12'h3b9;
			{5'd24, 5'd6}: color_data = 12'h3b9;
			{5'd24, 5'd7}: color_data = 12'h3b9;
			{5'd24, 5'd8}: color_data = 12'h752;
			{5'd24, 5'd9}: color_data = 12'h752;
			{5'd24, 5'd10}: color_data = 12'h752;
			{5'd24, 5'd11}: color_data = 12'h752;
			{5'd24, 5'd12}: color_data = 12'h752;
			{5'd24, 5'd13}: color_data = 12'h752;
			{5'd24, 5'd14}: color_data = 12'h752;
			{5'd24, 5'd15}: color_data = 12'h752;
			{5'd24, 5'd16}: color_data = 12'h752;
			{5'd24, 5'd17}: color_data = 12'h752;
			{5'd24, 5'd18}: color_data = 12'h852;
			{5'd24, 5'd19}: color_data = 12'h752;
			{5'd24, 5'd20}: color_data = 12'h3b9;
			{5'd24, 5'd21}: color_data = 12'h3b9;
			{5'd24, 5'd22}: color_data = 12'h000;
			{5'd24, 5'd23}: color_data = 12'h000;
			{5'd24, 5'd24}: color_data = 12'h000;
			{5'd24, 5'd25}: color_data = 12'h000;
			{5'd24, 5'd26}: color_data = 12'h000;
			{5'd24, 5'd27}: color_data = 12'h3b9;
			{5'd25, 5'd0}: color_data = 12'h3b9;
			{5'd25, 5'd1}: color_data = 12'h3b9;
			{5'd25, 5'd2}: color_data = 12'h3b9;
			{5'd25, 5'd3}: color_data = 12'h3b9;
			{5'd25, 5'd4}: color_data = 12'h3b9;
			{5'd25, 5'd5}: color_data = 12'h3b9;
			{5'd25, 5'd6}: color_data = 12'h3b9;
			{5'd25, 5'd7}: color_data = 12'h3b9;
			{5'd25, 5'd8}: color_data = 12'h752;
			{5'd25, 5'd9}: color_data = 12'h752;
			{5'd25, 5'd10}: color_data = 12'h752;
			{5'd25, 5'd11}: color_data = 12'h752;
			{5'd25, 5'd12}: color_data = 12'h752;
			{5'd25, 5'd13}: color_data = 12'h752;
			{5'd25, 5'd14}: color_data = 12'h752;
			{5'd25, 5'd15}: color_data = 12'h752;
			{5'd25, 5'd16}: color_data = 12'h752;
			{5'd25, 5'd17}: color_data = 12'h752;
			{5'd25, 5'd18}: color_data = 12'h752;
			{5'd25, 5'd19}: color_data = 12'h752;
			{5'd25, 5'd20}: color_data = 12'h3b9;
			{5'd25, 5'd21}: color_data = 12'h3b9;
			{5'd25, 5'd22}: color_data = 12'h000;
			{5'd25, 5'd23}: color_data = 12'h000;
			{5'd25, 5'd24}: color_data = 12'h000;
			{5'd25, 5'd25}: color_data = 12'h000;
			{5'd25, 5'd26}: color_data = 12'h000;
			{5'd25, 5'd27}: color_data = 12'h3b9;
			{5'd26, 5'd0}: color_data = 12'h3b9;
			{5'd26, 5'd1}: color_data = 12'h3b9;
			{5'd26, 5'd2}: color_data = 12'h3b9;
			{5'd26, 5'd3}: color_data = 12'h3b9;
			{5'd26, 5'd4}: color_data = 12'h3b9;
			{5'd26, 5'd5}: color_data = 12'h3b9;
			{5'd26, 5'd6}: color_data = 12'h3b9;
			{5'd26, 5'd7}: color_data = 12'h3b9;
			{5'd26, 5'd8}: color_data = 12'h3b9;
			{5'd26, 5'd9}: color_data = 12'h3b9;
			{5'd26, 5'd10}: color_data = 12'h3b9;
			{5'd26, 5'd11}: color_data = 12'h3b9;
			{5'd26, 5'd12}: color_data = 12'h752;
			{5'd26, 5'd13}: color_data = 12'h752;
			{5'd26, 5'd14}: color_data = 12'h752;
			{5'd26, 5'd15}: color_data = 12'h752;
			{5'd26, 5'd16}: color_data = 12'h752;
			{5'd26, 5'd17}: color_data = 12'h752;
			{5'd26, 5'd18}: color_data = 12'h3b9;
			{5'd26, 5'd19}: color_data = 12'h3b9;
			{5'd26, 5'd20}: color_data = 12'h3b9;
			{5'd26, 5'd21}: color_data = 12'h3b9;
			{5'd26, 5'd22}: color_data = 12'h3b9;
			{5'd26, 5'd23}: color_data = 12'h3b9;
			{5'd26, 5'd24}: color_data = 12'h3b9;
			{5'd26, 5'd25}: color_data = 12'h3b9;
			{5'd26, 5'd26}: color_data = 12'h3b9;
			{5'd26, 5'd27}: color_data = 12'h3b9;
            default: color_data = 12'h3b9;
        endcase
endmodule
