module intro_rom(
        input wire clk,
        input wire [7:0] x,
        input wire [7:0] y,
        output reg [11:0] color_data
);

    (* rom_style = "block" *)

    //signal declaration
    reg [7:0] x_reg;
    reg [7:0] y_reg;

    always @(posedge clk) begin
        x_reg <= x;
        y_reg <= y;
    end

    always @*
        case ({x_reg, y_reg})
			// right: 8'd171, bottom: 8'd159
			{8'd5, 8'd61}: color_data = 12'h000;
			{8'd5, 8'd62}: color_data = 12'h000;
			{8'd5, 8'd63}: color_data = 12'h000;
			{8'd5, 8'd64}: color_data = 12'h000;
			{8'd5, 8'd65}: color_data = 12'h000;
			{8'd5, 8'd66}: color_data = 12'h000;
			{8'd5, 8'd67}: color_data = 12'h000;
			{8'd5, 8'd68}: color_data = 12'h000;
			{8'd6, 8'd59}: color_data = 12'h000;
			{8'd6, 8'd60}: color_data = 12'h000;
			{8'd6, 8'd61}: color_data = 12'h000;
			{8'd6, 8'd62}: color_data = 12'h000;
			{8'd6, 8'd63}: color_data = 12'h000;
			{8'd6, 8'd64}: color_data = 12'h000;
			{8'd6, 8'd65}: color_data = 12'h000;
			{8'd6, 8'd66}: color_data = 12'h000;
			{8'd6, 8'd67}: color_data = 12'h000;
			{8'd6, 8'd68}: color_data = 12'h000;
			{8'd6, 8'd69}: color_data = 12'h000;
			{8'd7, 8'd56}: color_data = 12'h000;
			{8'd7, 8'd57}: color_data = 12'h000;
			{8'd7, 8'd58}: color_data = 12'h000;
			{8'd7, 8'd59}: color_data = 12'h000;
			{8'd7, 8'd60}: color_data = 12'h000;
			{8'd7, 8'd61}: color_data = 12'h000;
			{8'd7, 8'd62}: color_data = 12'h000;
			{8'd7, 8'd63}: color_data = 12'h000;
			{8'd7, 8'd64}: color_data = 12'h000;
			{8'd7, 8'd65}: color_data = 12'h000;
			{8'd7, 8'd66}: color_data = 12'h000;
			{8'd7, 8'd67}: color_data = 12'h000;
			{8'd7, 8'd68}: color_data = 12'h000;
			{8'd7, 8'd69}: color_data = 12'h000;
			{8'd8, 8'd54}: color_data = 12'h000;
			{8'd8, 8'd55}: color_data = 12'h000;
			{8'd8, 8'd56}: color_data = 12'h000;
			{8'd8, 8'd57}: color_data = 12'h000;
			{8'd8, 8'd58}: color_data = 12'h000;
			{8'd8, 8'd59}: color_data = 12'h000;
			{8'd8, 8'd60}: color_data = 12'h000;
			{8'd8, 8'd61}: color_data = 12'h200;
			{8'd8, 8'd62}: color_data = 12'h500;
			{8'd8, 8'd63}: color_data = 12'h000;
			{8'd8, 8'd64}: color_data = 12'h000;
			{8'd8, 8'd65}: color_data = 12'h000;
			{8'd8, 8'd66}: color_data = 12'h000;
			{8'd8, 8'd67}: color_data = 12'h000;
			{8'd8, 8'd68}: color_data = 12'h000;
			{8'd8, 8'd69}: color_data = 12'h000;
			{8'd8, 8'd70}: color_data = 12'h000;
			{8'd9, 8'd52}: color_data = 12'h000;
			{8'd9, 8'd53}: color_data = 12'h000;
			{8'd9, 8'd54}: color_data = 12'h000;
			{8'd9, 8'd55}: color_data = 12'h000;
			{8'd9, 8'd56}: color_data = 12'h000;
			{8'd9, 8'd57}: color_data = 12'h000;
			{8'd9, 8'd58}: color_data = 12'h000;
			{8'd9, 8'd59}: color_data = 12'h300;
			{8'd9, 8'd60}: color_data = 12'h910;
			{8'd9, 8'd61}: color_data = 12'hd20;
			{8'd9, 8'd62}: color_data = 12'hf21;
			{8'd9, 8'd63}: color_data = 12'h400;
			{8'd9, 8'd64}: color_data = 12'h000;
			{8'd9, 8'd65}: color_data = 12'h000;
			{8'd9, 8'd66}: color_data = 12'h000;
			{8'd9, 8'd67}: color_data = 12'h000;
			{8'd9, 8'd68}: color_data = 12'h000;
			{8'd9, 8'd69}: color_data = 12'h000;
			{8'd9, 8'd70}: color_data = 12'h000;
			{8'd10, 8'd49}: color_data = 12'h000;
			{8'd10, 8'd50}: color_data = 12'h000;
			{8'd10, 8'd51}: color_data = 12'h000;
			{8'd10, 8'd52}: color_data = 12'h000;
			{8'd10, 8'd53}: color_data = 12'h000;
			{8'd10, 8'd54}: color_data = 12'h000;
			{8'd10, 8'd55}: color_data = 12'h000;
			{8'd10, 8'd56}: color_data = 12'h000;
			{8'd10, 8'd57}: color_data = 12'h500;
			{8'd10, 8'd58}: color_data = 12'hb10;
			{8'd10, 8'd59}: color_data = 12'he21;
			{8'd10, 8'd60}: color_data = 12'he21;
			{8'd10, 8'd61}: color_data = 12'he21;
			{8'd10, 8'd62}: color_data = 12'he21;
			{8'd10, 8'd63}: color_data = 12'ha10;
			{8'd10, 8'd64}: color_data = 12'h000;
			{8'd10, 8'd65}: color_data = 12'h000;
			{8'd10, 8'd66}: color_data = 12'h000;
			{8'd10, 8'd67}: color_data = 12'h000;
			{8'd10, 8'd68}: color_data = 12'h000;
			{8'd10, 8'd69}: color_data = 12'h000;
			{8'd10, 8'd70}: color_data = 12'h000;
			{8'd11, 8'd47}: color_data = 12'h000;
			{8'd11, 8'd48}: color_data = 12'h000;
			{8'd11, 8'd49}: color_data = 12'h000;
			{8'd11, 8'd50}: color_data = 12'h000;
			{8'd11, 8'd51}: color_data = 12'h000;
			{8'd11, 8'd52}: color_data = 12'h000;
			{8'd11, 8'd53}: color_data = 12'h000;
			{8'd11, 8'd54}: color_data = 12'h200;
			{8'd11, 8'd55}: color_data = 12'h710;
			{8'd11, 8'd56}: color_data = 12'hc10;
			{8'd11, 8'd57}: color_data = 12'he21;
			{8'd11, 8'd58}: color_data = 12'he21;
			{8'd11, 8'd59}: color_data = 12'he21;
			{8'd11, 8'd60}: color_data = 12'he21;
			{8'd11, 8'd61}: color_data = 12'he21;
			{8'd11, 8'd62}: color_data = 12'he21;
			{8'd11, 8'd63}: color_data = 12'he21;
			{8'd11, 8'd64}: color_data = 12'h200;
			{8'd11, 8'd65}: color_data = 12'h000;
			{8'd11, 8'd66}: color_data = 12'h000;
			{8'd11, 8'd67}: color_data = 12'h000;
			{8'd11, 8'd68}: color_data = 12'h000;
			{8'd11, 8'd69}: color_data = 12'h000;
			{8'd11, 8'd70}: color_data = 12'h000;
			{8'd11, 8'd71}: color_data = 12'h000;
			{8'd11, 8'd120}: color_data = 12'hc00;
			{8'd11, 8'd121}: color_data = 12'hc01;
			{8'd11, 8'd122}: color_data = 12'hc01;
			{8'd11, 8'd123}: color_data = 12'he01;
			{8'd11, 8'd124}: color_data = 12'hb00;
			{8'd12, 8'd45}: color_data = 12'h000;
			{8'd12, 8'd46}: color_data = 12'h000;
			{8'd12, 8'd47}: color_data = 12'h000;
			{8'd12, 8'd48}: color_data = 12'h000;
			{8'd12, 8'd49}: color_data = 12'h000;
			{8'd12, 8'd50}: color_data = 12'h000;
			{8'd12, 8'd51}: color_data = 12'h000;
			{8'd12, 8'd52}: color_data = 12'h300;
			{8'd12, 8'd53}: color_data = 12'h910;
			{8'd12, 8'd54}: color_data = 12'hd20;
			{8'd12, 8'd55}: color_data = 12'he21;
			{8'd12, 8'd56}: color_data = 12'he21;
			{8'd12, 8'd57}: color_data = 12'he21;
			{8'd12, 8'd58}: color_data = 12'he21;
			{8'd12, 8'd59}: color_data = 12'he21;
			{8'd12, 8'd60}: color_data = 12'he21;
			{8'd12, 8'd61}: color_data = 12'he21;
			{8'd12, 8'd62}: color_data = 12'he21;
			{8'd12, 8'd63}: color_data = 12'he21;
			{8'd12, 8'd64}: color_data = 12'h810;
			{8'd12, 8'd65}: color_data = 12'h000;
			{8'd12, 8'd66}: color_data = 12'h000;
			{8'd12, 8'd67}: color_data = 12'h000;
			{8'd12, 8'd68}: color_data = 12'h000;
			{8'd12, 8'd69}: color_data = 12'h000;
			{8'd12, 8'd70}: color_data = 12'h000;
			{8'd12, 8'd71}: color_data = 12'h000;
			{8'd12, 8'd115}: color_data = 12'hc00;
			{8'd12, 8'd116}: color_data = 12'he00;
			{8'd12, 8'd117}: color_data = 12'he00;
			{8'd12, 8'd118}: color_data = 12'he00;
			{8'd12, 8'd119}: color_data = 12'he00;
			{8'd12, 8'd120}: color_data = 12'he00;
			{8'd12, 8'd121}: color_data = 12'he00;
			{8'd12, 8'd122}: color_data = 12'he00;
			{8'd12, 8'd123}: color_data = 12'he00;
			{8'd12, 8'd124}: color_data = 12'he00;
			{8'd12, 8'd125}: color_data = 12'he00;
			{8'd12, 8'd126}: color_data = 12'he00;
			{8'd12, 8'd127}: color_data = 12'he00;
			{8'd12, 8'd128}: color_data = 12'he00;
			{8'd12, 8'd129}: color_data = 12'hf00;
			{8'd13, 8'd42}: color_data = 12'h000;
			{8'd13, 8'd43}: color_data = 12'h000;
			{8'd13, 8'd44}: color_data = 12'h000;
			{8'd13, 8'd45}: color_data = 12'h000;
			{8'd13, 8'd46}: color_data = 12'h000;
			{8'd13, 8'd47}: color_data = 12'h000;
			{8'd13, 8'd48}: color_data = 12'h000;
			{8'd13, 8'd49}: color_data = 12'h000;
			{8'd13, 8'd50}: color_data = 12'h500;
			{8'd13, 8'd51}: color_data = 12'hb10;
			{8'd13, 8'd52}: color_data = 12'he21;
			{8'd13, 8'd53}: color_data = 12'he21;
			{8'd13, 8'd54}: color_data = 12'he21;
			{8'd13, 8'd55}: color_data = 12'he21;
			{8'd13, 8'd56}: color_data = 12'he21;
			{8'd13, 8'd57}: color_data = 12'he21;
			{8'd13, 8'd58}: color_data = 12'he21;
			{8'd13, 8'd59}: color_data = 12'he21;
			{8'd13, 8'd60}: color_data = 12'he21;
			{8'd13, 8'd61}: color_data = 12'he21;
			{8'd13, 8'd62}: color_data = 12'he21;
			{8'd13, 8'd63}: color_data = 12'he21;
			{8'd13, 8'd64}: color_data = 12'hd20;
			{8'd13, 8'd65}: color_data = 12'h100;
			{8'd13, 8'd66}: color_data = 12'h000;
			{8'd13, 8'd67}: color_data = 12'h000;
			{8'd13, 8'd68}: color_data = 12'h000;
			{8'd13, 8'd69}: color_data = 12'h000;
			{8'd13, 8'd70}: color_data = 12'h000;
			{8'd13, 8'd71}: color_data = 12'h000;
			{8'd13, 8'd72}: color_data = 12'h000;
			{8'd13, 8'd113}: color_data = 12'he01;
			{8'd13, 8'd114}: color_data = 12'he00;
			{8'd13, 8'd115}: color_data = 12'he00;
			{8'd13, 8'd116}: color_data = 12'he00;
			{8'd13, 8'd117}: color_data = 12'he01;
			{8'd13, 8'd118}: color_data = 12'he01;
			{8'd13, 8'd119}: color_data = 12'he00;
			{8'd13, 8'd120}: color_data = 12'he00;
			{8'd13, 8'd121}: color_data = 12'he00;
			{8'd13, 8'd122}: color_data = 12'he00;
			{8'd13, 8'd123}: color_data = 12'he00;
			{8'd13, 8'd124}: color_data = 12'he00;
			{8'd13, 8'd125}: color_data = 12'he01;
			{8'd13, 8'd126}: color_data = 12'he01;
			{8'd13, 8'd127}: color_data = 12'he00;
			{8'd13, 8'd128}: color_data = 12'he00;
			{8'd13, 8'd129}: color_data = 12'he00;
			{8'd13, 8'd130}: color_data = 12'he00;
			{8'd13, 8'd131}: color_data = 12'he00;
			{8'd14, 8'd40}: color_data = 12'h000;
			{8'd14, 8'd41}: color_data = 12'h000;
			{8'd14, 8'd42}: color_data = 12'h000;
			{8'd14, 8'd43}: color_data = 12'h000;
			{8'd14, 8'd44}: color_data = 12'h000;
			{8'd14, 8'd45}: color_data = 12'h000;
			{8'd14, 8'd46}: color_data = 12'h000;
			{8'd14, 8'd47}: color_data = 12'h200;
			{8'd14, 8'd48}: color_data = 12'h710;
			{8'd14, 8'd49}: color_data = 12'hc10;
			{8'd14, 8'd50}: color_data = 12'he21;
			{8'd14, 8'd51}: color_data = 12'he21;
			{8'd14, 8'd52}: color_data = 12'he21;
			{8'd14, 8'd53}: color_data = 12'he21;
			{8'd14, 8'd54}: color_data = 12'he21;
			{8'd14, 8'd55}: color_data = 12'he21;
			{8'd14, 8'd56}: color_data = 12'he21;
			{8'd14, 8'd57}: color_data = 12'he21;
			{8'd14, 8'd58}: color_data = 12'he21;
			{8'd14, 8'd59}: color_data = 12'he21;
			{8'd14, 8'd60}: color_data = 12'he21;
			{8'd14, 8'd61}: color_data = 12'he21;
			{8'd14, 8'd62}: color_data = 12'he21;
			{8'd14, 8'd63}: color_data = 12'he21;
			{8'd14, 8'd64}: color_data = 12'he21;
			{8'd14, 8'd65}: color_data = 12'h600;
			{8'd14, 8'd66}: color_data = 12'h000;
			{8'd14, 8'd67}: color_data = 12'h000;
			{8'd14, 8'd68}: color_data = 12'h000;
			{8'd14, 8'd69}: color_data = 12'h000;
			{8'd14, 8'd70}: color_data = 12'h000;
			{8'd14, 8'd71}: color_data = 12'h000;
			{8'd14, 8'd72}: color_data = 12'h000;
			{8'd14, 8'd111}: color_data = 12'he01;
			{8'd14, 8'd112}: color_data = 12'he00;
			{8'd14, 8'd113}: color_data = 12'he00;
			{8'd14, 8'd114}: color_data = 12'hf01;
			{8'd14, 8'd115}: color_data = 12'he00;
			{8'd14, 8'd116}: color_data = 12'he00;
			{8'd14, 8'd117}: color_data = 12'he00;
			{8'd14, 8'd118}: color_data = 12'he00;
			{8'd14, 8'd119}: color_data = 12'he00;
			{8'd14, 8'd120}: color_data = 12'he00;
			{8'd14, 8'd121}: color_data = 12'he00;
			{8'd14, 8'd122}: color_data = 12'he00;
			{8'd14, 8'd123}: color_data = 12'he00;
			{8'd14, 8'd124}: color_data = 12'he00;
			{8'd14, 8'd125}: color_data = 12'he00;
			{8'd14, 8'd126}: color_data = 12'he00;
			{8'd14, 8'd127}: color_data = 12'he00;
			{8'd14, 8'd128}: color_data = 12'he00;
			{8'd14, 8'd129}: color_data = 12'he00;
			{8'd14, 8'd130}: color_data = 12'he01;
			{8'd14, 8'd131}: color_data = 12'he00;
			{8'd14, 8'd132}: color_data = 12'he00;
			{8'd14, 8'd133}: color_data = 12'he00;
			{8'd15, 8'd38}: color_data = 12'h000;
			{8'd15, 8'd39}: color_data = 12'h000;
			{8'd15, 8'd40}: color_data = 12'h000;
			{8'd15, 8'd41}: color_data = 12'h000;
			{8'd15, 8'd42}: color_data = 12'h000;
			{8'd15, 8'd43}: color_data = 12'h000;
			{8'd15, 8'd44}: color_data = 12'h000;
			{8'd15, 8'd45}: color_data = 12'h300;
			{8'd15, 8'd46}: color_data = 12'h910;
			{8'd15, 8'd47}: color_data = 12'hd20;
			{8'd15, 8'd48}: color_data = 12'he21;
			{8'd15, 8'd49}: color_data = 12'he21;
			{8'd15, 8'd50}: color_data = 12'he21;
			{8'd15, 8'd51}: color_data = 12'he21;
			{8'd15, 8'd52}: color_data = 12'he21;
			{8'd15, 8'd53}: color_data = 12'he21;
			{8'd15, 8'd54}: color_data = 12'he21;
			{8'd15, 8'd55}: color_data = 12'he21;
			{8'd15, 8'd56}: color_data = 12'he21;
			{8'd15, 8'd57}: color_data = 12'he21;
			{8'd15, 8'd58}: color_data = 12'he21;
			{8'd15, 8'd59}: color_data = 12'he21;
			{8'd15, 8'd60}: color_data = 12'he21;
			{8'd15, 8'd61}: color_data = 12'he21;
			{8'd15, 8'd62}: color_data = 12'he21;
			{8'd15, 8'd63}: color_data = 12'he21;
			{8'd15, 8'd64}: color_data = 12'he21;
			{8'd15, 8'd65}: color_data = 12'hb10;
			{8'd15, 8'd66}: color_data = 12'h000;
			{8'd15, 8'd67}: color_data = 12'h000;
			{8'd15, 8'd68}: color_data = 12'h000;
			{8'd15, 8'd69}: color_data = 12'h000;
			{8'd15, 8'd70}: color_data = 12'h000;
			{8'd15, 8'd71}: color_data = 12'h000;
			{8'd15, 8'd72}: color_data = 12'h000;
			{8'd15, 8'd73}: color_data = 12'h000;
			{8'd15, 8'd109}: color_data = 12'hc00;
			{8'd15, 8'd110}: color_data = 12'he00;
			{8'd15, 8'd111}: color_data = 12'he00;
			{8'd15, 8'd112}: color_data = 12'hf01;
			{8'd15, 8'd113}: color_data = 12'he00;
			{8'd15, 8'd114}: color_data = 12'he00;
			{8'd15, 8'd115}: color_data = 12'he00;
			{8'd15, 8'd116}: color_data = 12'he00;
			{8'd15, 8'd117}: color_data = 12'he00;
			{8'd15, 8'd118}: color_data = 12'he00;
			{8'd15, 8'd119}: color_data = 12'he00;
			{8'd15, 8'd120}: color_data = 12'he00;
			{8'd15, 8'd121}: color_data = 12'he00;
			{8'd15, 8'd122}: color_data = 12'he00;
			{8'd15, 8'd123}: color_data = 12'he00;
			{8'd15, 8'd124}: color_data = 12'he00;
			{8'd15, 8'd125}: color_data = 12'he00;
			{8'd15, 8'd126}: color_data = 12'he00;
			{8'd15, 8'd127}: color_data = 12'he00;
			{8'd15, 8'd128}: color_data = 12'he00;
			{8'd15, 8'd129}: color_data = 12'he00;
			{8'd15, 8'd130}: color_data = 12'he00;
			{8'd15, 8'd131}: color_data = 12'he00;
			{8'd15, 8'd132}: color_data = 12'hf01;
			{8'd15, 8'd133}: color_data = 12'he00;
			{8'd15, 8'd134}: color_data = 12'he00;
			{8'd16, 8'd35}: color_data = 12'h000;
			{8'd16, 8'd36}: color_data = 12'h000;
			{8'd16, 8'd37}: color_data = 12'h000;
			{8'd16, 8'd38}: color_data = 12'h000;
			{8'd16, 8'd39}: color_data = 12'h000;
			{8'd16, 8'd40}: color_data = 12'h000;
			{8'd16, 8'd41}: color_data = 12'h000;
			{8'd16, 8'd42}: color_data = 12'h100;
			{8'd16, 8'd43}: color_data = 12'h500;
			{8'd16, 8'd44}: color_data = 12'hb10;
			{8'd16, 8'd45}: color_data = 12'he21;
			{8'd16, 8'd46}: color_data = 12'he21;
			{8'd16, 8'd47}: color_data = 12'he21;
			{8'd16, 8'd48}: color_data = 12'he21;
			{8'd16, 8'd49}: color_data = 12'he21;
			{8'd16, 8'd50}: color_data = 12'he21;
			{8'd16, 8'd51}: color_data = 12'he21;
			{8'd16, 8'd52}: color_data = 12'he21;
			{8'd16, 8'd53}: color_data = 12'he21;
			{8'd16, 8'd54}: color_data = 12'he21;
			{8'd16, 8'd55}: color_data = 12'he21;
			{8'd16, 8'd56}: color_data = 12'he21;
			{8'd16, 8'd57}: color_data = 12'he21;
			{8'd16, 8'd58}: color_data = 12'he21;
			{8'd16, 8'd59}: color_data = 12'he21;
			{8'd16, 8'd60}: color_data = 12'he21;
			{8'd16, 8'd61}: color_data = 12'he21;
			{8'd16, 8'd62}: color_data = 12'he21;
			{8'd16, 8'd63}: color_data = 12'he21;
			{8'd16, 8'd64}: color_data = 12'he21;
			{8'd16, 8'd65}: color_data = 12'he21;
			{8'd16, 8'd66}: color_data = 12'h400;
			{8'd16, 8'd67}: color_data = 12'h000;
			{8'd16, 8'd68}: color_data = 12'h000;
			{8'd16, 8'd69}: color_data = 12'h000;
			{8'd16, 8'd70}: color_data = 12'h000;
			{8'd16, 8'd71}: color_data = 12'h000;
			{8'd16, 8'd72}: color_data = 12'h000;
			{8'd16, 8'd73}: color_data = 12'h000;
			{8'd16, 8'd108}: color_data = 12'he01;
			{8'd16, 8'd109}: color_data = 12'he00;
			{8'd16, 8'd110}: color_data = 12'he01;
			{8'd16, 8'd111}: color_data = 12'he00;
			{8'd16, 8'd112}: color_data = 12'he00;
			{8'd16, 8'd113}: color_data = 12'he00;
			{8'd16, 8'd114}: color_data = 12'he00;
			{8'd16, 8'd115}: color_data = 12'he00;
			{8'd16, 8'd116}: color_data = 12'he00;
			{8'd16, 8'd117}: color_data = 12'he00;
			{8'd16, 8'd118}: color_data = 12'he00;
			{8'd16, 8'd119}: color_data = 12'he00;
			{8'd16, 8'd120}: color_data = 12'he01;
			{8'd16, 8'd121}: color_data = 12'he01;
			{8'd16, 8'd122}: color_data = 12'hf01;
			{8'd16, 8'd123}: color_data = 12'he01;
			{8'd16, 8'd124}: color_data = 12'he01;
			{8'd16, 8'd125}: color_data = 12'he00;
			{8'd16, 8'd126}: color_data = 12'he00;
			{8'd16, 8'd127}: color_data = 12'he00;
			{8'd16, 8'd128}: color_data = 12'he00;
			{8'd16, 8'd129}: color_data = 12'he00;
			{8'd16, 8'd130}: color_data = 12'he00;
			{8'd16, 8'd131}: color_data = 12'he00;
			{8'd16, 8'd132}: color_data = 12'he00;
			{8'd16, 8'd133}: color_data = 12'he00;
			{8'd16, 8'd134}: color_data = 12'he00;
			{8'd16, 8'd135}: color_data = 12'he00;
			{8'd16, 8'd136}: color_data = 12'he01;
			{8'd17, 8'd33}: color_data = 12'h000;
			{8'd17, 8'd34}: color_data = 12'h000;
			{8'd17, 8'd35}: color_data = 12'h000;
			{8'd17, 8'd36}: color_data = 12'h000;
			{8'd17, 8'd37}: color_data = 12'h000;
			{8'd17, 8'd38}: color_data = 12'h000;
			{8'd17, 8'd39}: color_data = 12'h000;
			{8'd17, 8'd40}: color_data = 12'h200;
			{8'd17, 8'd41}: color_data = 12'h710;
			{8'd17, 8'd42}: color_data = 12'hc10;
			{8'd17, 8'd43}: color_data = 12'he21;
			{8'd17, 8'd44}: color_data = 12'he21;
			{8'd17, 8'd45}: color_data = 12'he21;
			{8'd17, 8'd46}: color_data = 12'he21;
			{8'd17, 8'd47}: color_data = 12'he21;
			{8'd17, 8'd48}: color_data = 12'he21;
			{8'd17, 8'd49}: color_data = 12'he21;
			{8'd17, 8'd50}: color_data = 12'he21;
			{8'd17, 8'd51}: color_data = 12'he21;
			{8'd17, 8'd52}: color_data = 12'he21;
			{8'd17, 8'd53}: color_data = 12'he21;
			{8'd17, 8'd54}: color_data = 12'he21;
			{8'd17, 8'd55}: color_data = 12'he21;
			{8'd17, 8'd56}: color_data = 12'he21;
			{8'd17, 8'd57}: color_data = 12'he21;
			{8'd17, 8'd58}: color_data = 12'he21;
			{8'd17, 8'd59}: color_data = 12'he21;
			{8'd17, 8'd60}: color_data = 12'he21;
			{8'd17, 8'd61}: color_data = 12'he21;
			{8'd17, 8'd62}: color_data = 12'he21;
			{8'd17, 8'd63}: color_data = 12'he21;
			{8'd17, 8'd64}: color_data = 12'he21;
			{8'd17, 8'd65}: color_data = 12'he21;
			{8'd17, 8'd66}: color_data = 12'h910;
			{8'd17, 8'd67}: color_data = 12'h000;
			{8'd17, 8'd68}: color_data = 12'h000;
			{8'd17, 8'd69}: color_data = 12'h000;
			{8'd17, 8'd70}: color_data = 12'h000;
			{8'd17, 8'd71}: color_data = 12'h000;
			{8'd17, 8'd72}: color_data = 12'h000;
			{8'd17, 8'd73}: color_data = 12'h000;
			{8'd17, 8'd107}: color_data = 12'he00;
			{8'd17, 8'd108}: color_data = 12'he00;
			{8'd17, 8'd109}: color_data = 12'hf01;
			{8'd17, 8'd110}: color_data = 12'he00;
			{8'd17, 8'd111}: color_data = 12'he00;
			{8'd17, 8'd112}: color_data = 12'he00;
			{8'd17, 8'd113}: color_data = 12'he00;
			{8'd17, 8'd114}: color_data = 12'he00;
			{8'd17, 8'd115}: color_data = 12'he00;
			{8'd17, 8'd116}: color_data = 12'he01;
			{8'd17, 8'd117}: color_data = 12'he00;
			{8'd17, 8'd118}: color_data = 12'he00;
			{8'd17, 8'd119}: color_data = 12'he00;
			{8'd17, 8'd120}: color_data = 12'he00;
			{8'd17, 8'd121}: color_data = 12'he00;
			{8'd17, 8'd122}: color_data = 12'he00;
			{8'd17, 8'd123}: color_data = 12'he00;
			{8'd17, 8'd124}: color_data = 12'he00;
			{8'd17, 8'd125}: color_data = 12'he00;
			{8'd17, 8'd126}: color_data = 12'he00;
			{8'd17, 8'd127}: color_data = 12'he00;
			{8'd17, 8'd128}: color_data = 12'he01;
			{8'd17, 8'd129}: color_data = 12'he00;
			{8'd17, 8'd130}: color_data = 12'he00;
			{8'd17, 8'd131}: color_data = 12'he00;
			{8'd17, 8'd132}: color_data = 12'he00;
			{8'd17, 8'd133}: color_data = 12'he00;
			{8'd17, 8'd134}: color_data = 12'he00;
			{8'd17, 8'd135}: color_data = 12'hf01;
			{8'd17, 8'd136}: color_data = 12'he00;
			{8'd17, 8'd137}: color_data = 12'he00;
			{8'd18, 8'd31}: color_data = 12'h000;
			{8'd18, 8'd32}: color_data = 12'h000;
			{8'd18, 8'd33}: color_data = 12'h000;
			{8'd18, 8'd34}: color_data = 12'h000;
			{8'd18, 8'd35}: color_data = 12'h000;
			{8'd18, 8'd36}: color_data = 12'h000;
			{8'd18, 8'd37}: color_data = 12'h000;
			{8'd18, 8'd38}: color_data = 12'h300;
			{8'd18, 8'd39}: color_data = 12'h910;
			{8'd18, 8'd40}: color_data = 12'hd21;
			{8'd18, 8'd41}: color_data = 12'hf21;
			{8'd18, 8'd42}: color_data = 12'he21;
			{8'd18, 8'd43}: color_data = 12'he21;
			{8'd18, 8'd44}: color_data = 12'he21;
			{8'd18, 8'd45}: color_data = 12'he21;
			{8'd18, 8'd46}: color_data = 12'he21;
			{8'd18, 8'd47}: color_data = 12'he21;
			{8'd18, 8'd48}: color_data = 12'he21;
			{8'd18, 8'd49}: color_data = 12'he21;
			{8'd18, 8'd50}: color_data = 12'he21;
			{8'd18, 8'd51}: color_data = 12'he21;
			{8'd18, 8'd52}: color_data = 12'he21;
			{8'd18, 8'd53}: color_data = 12'he21;
			{8'd18, 8'd54}: color_data = 12'he21;
			{8'd18, 8'd55}: color_data = 12'he21;
			{8'd18, 8'd56}: color_data = 12'he21;
			{8'd18, 8'd57}: color_data = 12'he21;
			{8'd18, 8'd58}: color_data = 12'he21;
			{8'd18, 8'd59}: color_data = 12'he21;
			{8'd18, 8'd60}: color_data = 12'he21;
			{8'd18, 8'd61}: color_data = 12'he21;
			{8'd18, 8'd62}: color_data = 12'he21;
			{8'd18, 8'd63}: color_data = 12'he21;
			{8'd18, 8'd64}: color_data = 12'he21;
			{8'd18, 8'd65}: color_data = 12'he21;
			{8'd18, 8'd66}: color_data = 12'hd20;
			{8'd18, 8'd67}: color_data = 12'h200;
			{8'd18, 8'd68}: color_data = 12'h000;
			{8'd18, 8'd69}: color_data = 12'h000;
			{8'd18, 8'd70}: color_data = 12'h000;
			{8'd18, 8'd71}: color_data = 12'h000;
			{8'd18, 8'd72}: color_data = 12'h000;
			{8'd18, 8'd73}: color_data = 12'h000;
			{8'd18, 8'd74}: color_data = 12'h000;
			{8'd18, 8'd106}: color_data = 12'he00;
			{8'd18, 8'd107}: color_data = 12'he00;
			{8'd18, 8'd108}: color_data = 12'he00;
			{8'd18, 8'd109}: color_data = 12'he00;
			{8'd18, 8'd110}: color_data = 12'he00;
			{8'd18, 8'd111}: color_data = 12'he00;
			{8'd18, 8'd112}: color_data = 12'he00;
			{8'd18, 8'd113}: color_data = 12'he00;
			{8'd18, 8'd114}: color_data = 12'he01;
			{8'd18, 8'd115}: color_data = 12'he00;
			{8'd18, 8'd116}: color_data = 12'he00;
			{8'd18, 8'd117}: color_data = 12'he00;
			{8'd18, 8'd118}: color_data = 12'he00;
			{8'd18, 8'd125}: color_data = 12'hf00;
			{8'd18, 8'd126}: color_data = 12'he00;
			{8'd18, 8'd127}: color_data = 12'he00;
			{8'd18, 8'd128}: color_data = 12'he00;
			{8'd18, 8'd129}: color_data = 12'he00;
			{8'd18, 8'd130}: color_data = 12'he01;
			{8'd18, 8'd131}: color_data = 12'he00;
			{8'd18, 8'd132}: color_data = 12'he00;
			{8'd18, 8'd133}: color_data = 12'he00;
			{8'd18, 8'd134}: color_data = 12'he00;
			{8'd18, 8'd135}: color_data = 12'he00;
			{8'd18, 8'd136}: color_data = 12'he01;
			{8'd18, 8'd137}: color_data = 12'he00;
			{8'd18, 8'd138}: color_data = 12'hd00;
			{8'd19, 8'd29}: color_data = 12'h000;
			{8'd19, 8'd30}: color_data = 12'h000;
			{8'd19, 8'd31}: color_data = 12'h000;
			{8'd19, 8'd32}: color_data = 12'h000;
			{8'd19, 8'd33}: color_data = 12'h000;
			{8'd19, 8'd34}: color_data = 12'h000;
			{8'd19, 8'd35}: color_data = 12'h100;
			{8'd19, 8'd36}: color_data = 12'h500;
			{8'd19, 8'd37}: color_data = 12'hb10;
			{8'd19, 8'd38}: color_data = 12'he21;
			{8'd19, 8'd39}: color_data = 12'he21;
			{8'd19, 8'd40}: color_data = 12'he21;
			{8'd19, 8'd41}: color_data = 12'he21;
			{8'd19, 8'd42}: color_data = 12'he21;
			{8'd19, 8'd43}: color_data = 12'he21;
			{8'd19, 8'd44}: color_data = 12'he21;
			{8'd19, 8'd45}: color_data = 12'he21;
			{8'd19, 8'd46}: color_data = 12'he21;
			{8'd19, 8'd47}: color_data = 12'he21;
			{8'd19, 8'd48}: color_data = 12'he21;
			{8'd19, 8'd49}: color_data = 12'he21;
			{8'd19, 8'd50}: color_data = 12'he21;
			{8'd19, 8'd51}: color_data = 12'he21;
			{8'd19, 8'd52}: color_data = 12'he21;
			{8'd19, 8'd53}: color_data = 12'he21;
			{8'd19, 8'd54}: color_data = 12'he21;
			{8'd19, 8'd55}: color_data = 12'he21;
			{8'd19, 8'd56}: color_data = 12'he21;
			{8'd19, 8'd57}: color_data = 12'he21;
			{8'd19, 8'd58}: color_data = 12'he21;
			{8'd19, 8'd59}: color_data = 12'he21;
			{8'd19, 8'd60}: color_data = 12'he21;
			{8'd19, 8'd61}: color_data = 12'he21;
			{8'd19, 8'd62}: color_data = 12'he21;
			{8'd19, 8'd63}: color_data = 12'he21;
			{8'd19, 8'd64}: color_data = 12'he21;
			{8'd19, 8'd65}: color_data = 12'he21;
			{8'd19, 8'd66}: color_data = 12'hf21;
			{8'd19, 8'd67}: color_data = 12'h810;
			{8'd19, 8'd68}: color_data = 12'h000;
			{8'd19, 8'd69}: color_data = 12'h000;
			{8'd19, 8'd70}: color_data = 12'h000;
			{8'd19, 8'd71}: color_data = 12'h000;
			{8'd19, 8'd72}: color_data = 12'h000;
			{8'd19, 8'd73}: color_data = 12'h000;
			{8'd19, 8'd74}: color_data = 12'h000;
			{8'd19, 8'd105}: color_data = 12'he00;
			{8'd19, 8'd106}: color_data = 12'he00;
			{8'd19, 8'd107}: color_data = 12'he00;
			{8'd19, 8'd108}: color_data = 12'he00;
			{8'd19, 8'd109}: color_data = 12'he00;
			{8'd19, 8'd110}: color_data = 12'he00;
			{8'd19, 8'd111}: color_data = 12'he00;
			{8'd19, 8'd112}: color_data = 12'he01;
			{8'd19, 8'd113}: color_data = 12'he00;
			{8'd19, 8'd114}: color_data = 12'he00;
			{8'd19, 8'd115}: color_data = 12'he01;
			{8'd19, 8'd129}: color_data = 12'he00;
			{8'd19, 8'd130}: color_data = 12'he00;
			{8'd19, 8'd131}: color_data = 12'he00;
			{8'd19, 8'd132}: color_data = 12'he00;
			{8'd19, 8'd133}: color_data = 12'he00;
			{8'd19, 8'd134}: color_data = 12'he00;
			{8'd19, 8'd135}: color_data = 12'he00;
			{8'd19, 8'd136}: color_data = 12'he00;
			{8'd19, 8'd137}: color_data = 12'he00;
			{8'd19, 8'd138}: color_data = 12'he00;
			{8'd19, 8'd139}: color_data = 12'hd00;
			{8'd20, 8'd29}: color_data = 12'h000;
			{8'd20, 8'd30}: color_data = 12'h000;
			{8'd20, 8'd31}: color_data = 12'h000;
			{8'd20, 8'd32}: color_data = 12'h000;
			{8'd20, 8'd33}: color_data = 12'h200;
			{8'd20, 8'd34}: color_data = 12'h710;
			{8'd20, 8'd35}: color_data = 12'hc10;
			{8'd20, 8'd36}: color_data = 12'he21;
			{8'd20, 8'd37}: color_data = 12'he21;
			{8'd20, 8'd38}: color_data = 12'he21;
			{8'd20, 8'd39}: color_data = 12'he21;
			{8'd20, 8'd40}: color_data = 12'he21;
			{8'd20, 8'd41}: color_data = 12'he21;
			{8'd20, 8'd42}: color_data = 12'he21;
			{8'd20, 8'd43}: color_data = 12'he21;
			{8'd20, 8'd44}: color_data = 12'he21;
			{8'd20, 8'd45}: color_data = 12'he21;
			{8'd20, 8'd46}: color_data = 12'he21;
			{8'd20, 8'd47}: color_data = 12'he21;
			{8'd20, 8'd48}: color_data = 12'he21;
			{8'd20, 8'd49}: color_data = 12'he21;
			{8'd20, 8'd50}: color_data = 12'he21;
			{8'd20, 8'd51}: color_data = 12'he21;
			{8'd20, 8'd52}: color_data = 12'he21;
			{8'd20, 8'd53}: color_data = 12'he21;
			{8'd20, 8'd54}: color_data = 12'he21;
			{8'd20, 8'd55}: color_data = 12'he21;
			{8'd20, 8'd56}: color_data = 12'he21;
			{8'd20, 8'd57}: color_data = 12'he21;
			{8'd20, 8'd58}: color_data = 12'he21;
			{8'd20, 8'd59}: color_data = 12'he21;
			{8'd20, 8'd60}: color_data = 12'he21;
			{8'd20, 8'd61}: color_data = 12'he21;
			{8'd20, 8'd62}: color_data = 12'he21;
			{8'd20, 8'd63}: color_data = 12'he21;
			{8'd20, 8'd64}: color_data = 12'he21;
			{8'd20, 8'd65}: color_data = 12'he21;
			{8'd20, 8'd66}: color_data = 12'hd20;
			{8'd20, 8'd67}: color_data = 12'h810;
			{8'd20, 8'd68}: color_data = 12'h000;
			{8'd20, 8'd69}: color_data = 12'h000;
			{8'd20, 8'd70}: color_data = 12'h000;
			{8'd20, 8'd71}: color_data = 12'h000;
			{8'd20, 8'd72}: color_data = 12'h000;
			{8'd20, 8'd73}: color_data = 12'h000;
			{8'd20, 8'd74}: color_data = 12'h000;
			{8'd20, 8'd75}: color_data = 12'h000;
			{8'd20, 8'd104}: color_data = 12'hd00;
			{8'd20, 8'd105}: color_data = 12'he00;
			{8'd20, 8'd106}: color_data = 12'he00;
			{8'd20, 8'd107}: color_data = 12'he00;
			{8'd20, 8'd108}: color_data = 12'he00;
			{8'd20, 8'd109}: color_data = 12'he00;
			{8'd20, 8'd110}: color_data = 12'he00;
			{8'd20, 8'd111}: color_data = 12'he01;
			{8'd20, 8'd112}: color_data = 12'he00;
			{8'd20, 8'd113}: color_data = 12'he01;
			{8'd20, 8'd131}: color_data = 12'he01;
			{8'd20, 8'd132}: color_data = 12'he00;
			{8'd20, 8'd133}: color_data = 12'he01;
			{8'd20, 8'd134}: color_data = 12'he00;
			{8'd20, 8'd135}: color_data = 12'he00;
			{8'd20, 8'd136}: color_data = 12'he00;
			{8'd20, 8'd137}: color_data = 12'he00;
			{8'd20, 8'd138}: color_data = 12'hf01;
			{8'd20, 8'd139}: color_data = 12'he00;
			{8'd20, 8'd140}: color_data = 12'hf00;
			{8'd21, 8'd30}: color_data = 12'h000;
			{8'd21, 8'd31}: color_data = 12'h000;
			{8'd21, 8'd32}: color_data = 12'h100;
			{8'd21, 8'd33}: color_data = 12'hd20;
			{8'd21, 8'd34}: color_data = 12'hf21;
			{8'd21, 8'd35}: color_data = 12'he21;
			{8'd21, 8'd36}: color_data = 12'he21;
			{8'd21, 8'd37}: color_data = 12'he21;
			{8'd21, 8'd38}: color_data = 12'he21;
			{8'd21, 8'd39}: color_data = 12'he21;
			{8'd21, 8'd40}: color_data = 12'he21;
			{8'd21, 8'd41}: color_data = 12'he21;
			{8'd21, 8'd42}: color_data = 12'he21;
			{8'd21, 8'd43}: color_data = 12'he21;
			{8'd21, 8'd44}: color_data = 12'he21;
			{8'd21, 8'd45}: color_data = 12'he21;
			{8'd21, 8'd46}: color_data = 12'he21;
			{8'd21, 8'd47}: color_data = 12'he21;
			{8'd21, 8'd48}: color_data = 12'he21;
			{8'd21, 8'd49}: color_data = 12'he21;
			{8'd21, 8'd50}: color_data = 12'he21;
			{8'd21, 8'd51}: color_data = 12'he21;
			{8'd21, 8'd52}: color_data = 12'he21;
			{8'd21, 8'd53}: color_data = 12'he21;
			{8'd21, 8'd54}: color_data = 12'he21;
			{8'd21, 8'd55}: color_data = 12'he21;
			{8'd21, 8'd56}: color_data = 12'he21;
			{8'd21, 8'd57}: color_data = 12'he21;
			{8'd21, 8'd58}: color_data = 12'he21;
			{8'd21, 8'd59}: color_data = 12'he21;
			{8'd21, 8'd60}: color_data = 12'he21;
			{8'd21, 8'd61}: color_data = 12'he21;
			{8'd21, 8'd62}: color_data = 12'he21;
			{8'd21, 8'd63}: color_data = 12'hd20;
			{8'd21, 8'd64}: color_data = 12'h910;
			{8'd21, 8'd65}: color_data = 12'h500;
			{8'd21, 8'd66}: color_data = 12'h100;
			{8'd21, 8'd67}: color_data = 12'h000;
			{8'd21, 8'd68}: color_data = 12'h000;
			{8'd21, 8'd69}: color_data = 12'h000;
			{8'd21, 8'd70}: color_data = 12'h000;
			{8'd21, 8'd71}: color_data = 12'h000;
			{8'd21, 8'd72}: color_data = 12'h000;
			{8'd21, 8'd73}: color_data = 12'h000;
			{8'd21, 8'd74}: color_data = 12'h000;
			{8'd21, 8'd75}: color_data = 12'h000;
			{8'd21, 8'd104}: color_data = 12'he00;
			{8'd21, 8'd105}: color_data = 12'hf00;
			{8'd21, 8'd106}: color_data = 12'he00;
			{8'd21, 8'd107}: color_data = 12'he00;
			{8'd21, 8'd108}: color_data = 12'he00;
			{8'd21, 8'd109}: color_data = 12'he00;
			{8'd21, 8'd110}: color_data = 12'he01;
			{8'd21, 8'd111}: color_data = 12'he00;
			{8'd21, 8'd112}: color_data = 12'he01;
			{8'd21, 8'd132}: color_data = 12'hd00;
			{8'd21, 8'd133}: color_data = 12'he00;
			{8'd21, 8'd134}: color_data = 12'he01;
			{8'd21, 8'd135}: color_data = 12'he00;
			{8'd21, 8'd136}: color_data = 12'he00;
			{8'd21, 8'd137}: color_data = 12'he00;
			{8'd21, 8'd138}: color_data = 12'he00;
			{8'd21, 8'd139}: color_data = 12'he00;
			{8'd21, 8'd140}: color_data = 12'he00;
			{8'd22, 8'd30}: color_data = 12'h000;
			{8'd22, 8'd31}: color_data = 12'h000;
			{8'd22, 8'd32}: color_data = 12'h100;
			{8'd22, 8'd33}: color_data = 12'hd20;
			{8'd22, 8'd34}: color_data = 12'he21;
			{8'd22, 8'd35}: color_data = 12'he21;
			{8'd22, 8'd36}: color_data = 12'he21;
			{8'd22, 8'd37}: color_data = 12'he21;
			{8'd22, 8'd38}: color_data = 12'he21;
			{8'd22, 8'd39}: color_data = 12'he21;
			{8'd22, 8'd40}: color_data = 12'he21;
			{8'd22, 8'd41}: color_data = 12'he21;
			{8'd22, 8'd42}: color_data = 12'he21;
			{8'd22, 8'd43}: color_data = 12'he21;
			{8'd22, 8'd44}: color_data = 12'he21;
			{8'd22, 8'd45}: color_data = 12'he21;
			{8'd22, 8'd46}: color_data = 12'he21;
			{8'd22, 8'd47}: color_data = 12'he21;
			{8'd22, 8'd48}: color_data = 12'he21;
			{8'd22, 8'd49}: color_data = 12'he21;
			{8'd22, 8'd50}: color_data = 12'he21;
			{8'd22, 8'd51}: color_data = 12'he21;
			{8'd22, 8'd52}: color_data = 12'he21;
			{8'd22, 8'd53}: color_data = 12'he21;
			{8'd22, 8'd54}: color_data = 12'he21;
			{8'd22, 8'd55}: color_data = 12'he21;
			{8'd22, 8'd56}: color_data = 12'he21;
			{8'd22, 8'd57}: color_data = 12'he21;
			{8'd22, 8'd58}: color_data = 12'he21;
			{8'd22, 8'd59}: color_data = 12'he21;
			{8'd22, 8'd60}: color_data = 12'hc10;
			{8'd22, 8'd61}: color_data = 12'h810;
			{8'd22, 8'd62}: color_data = 12'h400;
			{8'd22, 8'd63}: color_data = 12'h100;
			{8'd22, 8'd64}: color_data = 12'h000;
			{8'd22, 8'd65}: color_data = 12'h000;
			{8'd22, 8'd66}: color_data = 12'h000;
			{8'd22, 8'd67}: color_data = 12'h000;
			{8'd22, 8'd68}: color_data = 12'h000;
			{8'd22, 8'd69}: color_data = 12'h000;
			{8'd22, 8'd70}: color_data = 12'h000;
			{8'd22, 8'd71}: color_data = 12'h000;
			{8'd22, 8'd72}: color_data = 12'h000;
			{8'd22, 8'd73}: color_data = 12'h000;
			{8'd22, 8'd74}: color_data = 12'h000;
			{8'd22, 8'd75}: color_data = 12'h000;
			{8'd22, 8'd103}: color_data = 12'he00;
			{8'd22, 8'd104}: color_data = 12'he00;
			{8'd22, 8'd105}: color_data = 12'he00;
			{8'd22, 8'd106}: color_data = 12'he00;
			{8'd22, 8'd107}: color_data = 12'he00;
			{8'd22, 8'd108}: color_data = 12'he00;
			{8'd22, 8'd109}: color_data = 12'he00;
			{8'd22, 8'd110}: color_data = 12'he00;
			{8'd22, 8'd111}: color_data = 12'hf00;
			{8'd22, 8'd133}: color_data = 12'he01;
			{8'd22, 8'd134}: color_data = 12'he00;
			{8'd22, 8'd135}: color_data = 12'he00;
			{8'd22, 8'd136}: color_data = 12'he00;
			{8'd22, 8'd137}: color_data = 12'he00;
			{8'd22, 8'd138}: color_data = 12'he00;
			{8'd22, 8'd139}: color_data = 12'he00;
			{8'd22, 8'd140}: color_data = 12'he00;
			{8'd22, 8'd141}: color_data = 12'he01;
			{8'd23, 8'd30}: color_data = 12'h000;
			{8'd23, 8'd31}: color_data = 12'h000;
			{8'd23, 8'd32}: color_data = 12'h000;
			{8'd23, 8'd33}: color_data = 12'hb10;
			{8'd23, 8'd34}: color_data = 12'he21;
			{8'd23, 8'd35}: color_data = 12'he21;
			{8'd23, 8'd36}: color_data = 12'he21;
			{8'd23, 8'd37}: color_data = 12'he21;
			{8'd23, 8'd38}: color_data = 12'he21;
			{8'd23, 8'd39}: color_data = 12'he21;
			{8'd23, 8'd40}: color_data = 12'he21;
			{8'd23, 8'd41}: color_data = 12'he21;
			{8'd23, 8'd42}: color_data = 12'he21;
			{8'd23, 8'd43}: color_data = 12'he21;
			{8'd23, 8'd44}: color_data = 12'he21;
			{8'd23, 8'd45}: color_data = 12'he21;
			{8'd23, 8'd46}: color_data = 12'he21;
			{8'd23, 8'd47}: color_data = 12'he21;
			{8'd23, 8'd48}: color_data = 12'he21;
			{8'd23, 8'd49}: color_data = 12'he21;
			{8'd23, 8'd50}: color_data = 12'he21;
			{8'd23, 8'd51}: color_data = 12'he21;
			{8'd23, 8'd52}: color_data = 12'he21;
			{8'd23, 8'd53}: color_data = 12'he21;
			{8'd23, 8'd54}: color_data = 12'he21;
			{8'd23, 8'd55}: color_data = 12'he21;
			{8'd23, 8'd56}: color_data = 12'he20;
			{8'd23, 8'd57}: color_data = 12'hb10;
			{8'd23, 8'd58}: color_data = 12'h710;
			{8'd23, 8'd59}: color_data = 12'h300;
			{8'd23, 8'd60}: color_data = 12'h000;
			{8'd23, 8'd61}: color_data = 12'h000;
			{8'd23, 8'd62}: color_data = 12'h000;
			{8'd23, 8'd63}: color_data = 12'h000;
			{8'd23, 8'd64}: color_data = 12'h000;
			{8'd23, 8'd65}: color_data = 12'h000;
			{8'd23, 8'd66}: color_data = 12'h000;
			{8'd23, 8'd67}: color_data = 12'h000;
			{8'd23, 8'd68}: color_data = 12'h000;
			{8'd23, 8'd69}: color_data = 12'h000;
			{8'd23, 8'd70}: color_data = 12'h000;
			{8'd23, 8'd71}: color_data = 12'h000;
			{8'd23, 8'd72}: color_data = 12'h000;
			{8'd23, 8'd73}: color_data = 12'h000;
			{8'd23, 8'd102}: color_data = 12'hd01;
			{8'd23, 8'd103}: color_data = 12'he00;
			{8'd23, 8'd104}: color_data = 12'he00;
			{8'd23, 8'd105}: color_data = 12'he00;
			{8'd23, 8'd106}: color_data = 12'he00;
			{8'd23, 8'd107}: color_data = 12'he00;
			{8'd23, 8'd108}: color_data = 12'he01;
			{8'd23, 8'd109}: color_data = 12'he00;
			{8'd23, 8'd110}: color_data = 12'hf00;
			{8'd23, 8'd134}: color_data = 12'hd01;
			{8'd23, 8'd135}: color_data = 12'he00;
			{8'd23, 8'd136}: color_data = 12'he00;
			{8'd23, 8'd137}: color_data = 12'he00;
			{8'd23, 8'd138}: color_data = 12'he00;
			{8'd23, 8'd139}: color_data = 12'he00;
			{8'd23, 8'd140}: color_data = 12'he00;
			{8'd23, 8'd141}: color_data = 12'he00;
			{8'd24, 8'd22}: color_data = 12'h000;
			{8'd24, 8'd23}: color_data = 12'h000;
			{8'd24, 8'd24}: color_data = 12'h000;
			{8'd24, 8'd25}: color_data = 12'h000;
			{8'd24, 8'd26}: color_data = 12'h000;
			{8'd24, 8'd27}: color_data = 12'h000;
			{8'd24, 8'd28}: color_data = 12'h000;
			{8'd24, 8'd30}: color_data = 12'h000;
			{8'd24, 8'd31}: color_data = 12'h000;
			{8'd24, 8'd32}: color_data = 12'h000;
			{8'd24, 8'd33}: color_data = 12'ha10;
			{8'd24, 8'd34}: color_data = 12'he21;
			{8'd24, 8'd35}: color_data = 12'he21;
			{8'd24, 8'd36}: color_data = 12'he21;
			{8'd24, 8'd37}: color_data = 12'he21;
			{8'd24, 8'd38}: color_data = 12'he21;
			{8'd24, 8'd39}: color_data = 12'he21;
			{8'd24, 8'd40}: color_data = 12'he21;
			{8'd24, 8'd41}: color_data = 12'he21;
			{8'd24, 8'd42}: color_data = 12'he21;
			{8'd24, 8'd43}: color_data = 12'he21;
			{8'd24, 8'd44}: color_data = 12'he21;
			{8'd24, 8'd45}: color_data = 12'he21;
			{8'd24, 8'd46}: color_data = 12'he21;
			{8'd24, 8'd47}: color_data = 12'he21;
			{8'd24, 8'd48}: color_data = 12'he21;
			{8'd24, 8'd49}: color_data = 12'he21;
			{8'd24, 8'd50}: color_data = 12'he21;
			{8'd24, 8'd51}: color_data = 12'he21;
			{8'd24, 8'd52}: color_data = 12'he21;
			{8'd24, 8'd53}: color_data = 12'hd20;
			{8'd24, 8'd54}: color_data = 12'ha10;
			{8'd24, 8'd55}: color_data = 12'h600;
			{8'd24, 8'd56}: color_data = 12'h200;
			{8'd24, 8'd57}: color_data = 12'h000;
			{8'd24, 8'd58}: color_data = 12'h000;
			{8'd24, 8'd59}: color_data = 12'h000;
			{8'd24, 8'd60}: color_data = 12'h000;
			{8'd24, 8'd61}: color_data = 12'h000;
			{8'd24, 8'd62}: color_data = 12'h000;
			{8'd24, 8'd63}: color_data = 12'h000;
			{8'd24, 8'd64}: color_data = 12'h000;
			{8'd24, 8'd65}: color_data = 12'h000;
			{8'd24, 8'd66}: color_data = 12'h000;
			{8'd24, 8'd67}: color_data = 12'h000;
			{8'd24, 8'd68}: color_data = 12'h000;
			{8'd24, 8'd69}: color_data = 12'h000;
			{8'd24, 8'd70}: color_data = 12'h000;
			{8'd24, 8'd102}: color_data = 12'he00;
			{8'd24, 8'd103}: color_data = 12'he00;
			{8'd24, 8'd104}: color_data = 12'he00;
			{8'd24, 8'd105}: color_data = 12'he00;
			{8'd24, 8'd106}: color_data = 12'he00;
			{8'd24, 8'd107}: color_data = 12'he00;
			{8'd24, 8'd108}: color_data = 12'he00;
			{8'd24, 8'd109}: color_data = 12'he00;
			{8'd24, 8'd135}: color_data = 12'he00;
			{8'd24, 8'd136}: color_data = 12'he00;
			{8'd24, 8'd137}: color_data = 12'he00;
			{8'd24, 8'd138}: color_data = 12'he00;
			{8'd24, 8'd139}: color_data = 12'he00;
			{8'd24, 8'd140}: color_data = 12'he00;
			{8'd24, 8'd141}: color_data = 12'he00;
			{8'd24, 8'd142}: color_data = 12'he01;
			{8'd25, 8'd11}: color_data = 12'h000;
			{8'd25, 8'd12}: color_data = 12'h000;
			{8'd25, 8'd13}: color_data = 12'h000;
			{8'd25, 8'd14}: color_data = 12'h000;
			{8'd25, 8'd15}: color_data = 12'h000;
			{8'd25, 8'd16}: color_data = 12'h000;
			{8'd25, 8'd21}: color_data = 12'h000;
			{8'd25, 8'd22}: color_data = 12'h000;
			{8'd25, 8'd23}: color_data = 12'h000;
			{8'd25, 8'd24}: color_data = 12'h000;
			{8'd25, 8'd25}: color_data = 12'h000;
			{8'd25, 8'd26}: color_data = 12'h000;
			{8'd25, 8'd27}: color_data = 12'h000;
			{8'd25, 8'd28}: color_data = 12'h000;
			{8'd25, 8'd30}: color_data = 12'h000;
			{8'd25, 8'd31}: color_data = 12'h000;
			{8'd25, 8'd32}: color_data = 12'h000;
			{8'd25, 8'd33}: color_data = 12'h810;
			{8'd25, 8'd34}: color_data = 12'he21;
			{8'd25, 8'd35}: color_data = 12'he21;
			{8'd25, 8'd36}: color_data = 12'he21;
			{8'd25, 8'd37}: color_data = 12'he21;
			{8'd25, 8'd38}: color_data = 12'he21;
			{8'd25, 8'd39}: color_data = 12'he21;
			{8'd25, 8'd40}: color_data = 12'he21;
			{8'd25, 8'd41}: color_data = 12'he21;
			{8'd25, 8'd42}: color_data = 12'he21;
			{8'd25, 8'd43}: color_data = 12'he21;
			{8'd25, 8'd44}: color_data = 12'he21;
			{8'd25, 8'd45}: color_data = 12'he21;
			{8'd25, 8'd46}: color_data = 12'he21;
			{8'd25, 8'd47}: color_data = 12'he21;
			{8'd25, 8'd48}: color_data = 12'he21;
			{8'd25, 8'd49}: color_data = 12'he21;
			{8'd25, 8'd50}: color_data = 12'hc10;
			{8'd25, 8'd51}: color_data = 12'h910;
			{8'd25, 8'd52}: color_data = 12'h500;
			{8'd25, 8'd53}: color_data = 12'h100;
			{8'd25, 8'd54}: color_data = 12'h000;
			{8'd25, 8'd55}: color_data = 12'h000;
			{8'd25, 8'd56}: color_data = 12'h000;
			{8'd25, 8'd57}: color_data = 12'h000;
			{8'd25, 8'd58}: color_data = 12'h000;
			{8'd25, 8'd59}: color_data = 12'h000;
			{8'd25, 8'd60}: color_data = 12'h000;
			{8'd25, 8'd61}: color_data = 12'h000;
			{8'd25, 8'd62}: color_data = 12'h000;
			{8'd25, 8'd63}: color_data = 12'h000;
			{8'd25, 8'd64}: color_data = 12'h000;
			{8'd25, 8'd65}: color_data = 12'h000;
			{8'd25, 8'd66}: color_data = 12'h000;
			{8'd25, 8'd67}: color_data = 12'h000;
			{8'd25, 8'd101}: color_data = 12'hc00;
			{8'd25, 8'd102}: color_data = 12'he00;
			{8'd25, 8'd103}: color_data = 12'he00;
			{8'd25, 8'd104}: color_data = 12'he00;
			{8'd25, 8'd105}: color_data = 12'he00;
			{8'd25, 8'd106}: color_data = 12'he00;
			{8'd25, 8'd107}: color_data = 12'he00;
			{8'd25, 8'd108}: color_data = 12'he00;
			{8'd25, 8'd136}: color_data = 12'he01;
			{8'd25, 8'd137}: color_data = 12'he01;
			{8'd25, 8'd138}: color_data = 12'he00;
			{8'd25, 8'd139}: color_data = 12'he00;
			{8'd25, 8'd140}: color_data = 12'he00;
			{8'd25, 8'd141}: color_data = 12'he01;
			{8'd25, 8'd142}: color_data = 12'he00;
			{8'd26, 8'd10}: color_data = 12'h000;
			{8'd26, 8'd11}: color_data = 12'h000;
			{8'd26, 8'd12}: color_data = 12'h000;
			{8'd26, 8'd13}: color_data = 12'h000;
			{8'd26, 8'd14}: color_data = 12'h000;
			{8'd26, 8'd15}: color_data = 12'h000;
			{8'd26, 8'd16}: color_data = 12'h000;
			{8'd26, 8'd17}: color_data = 12'h000;
			{8'd26, 8'd20}: color_data = 12'h000;
			{8'd26, 8'd21}: color_data = 12'h000;
			{8'd26, 8'd22}: color_data = 12'h000;
			{8'd26, 8'd23}: color_data = 12'h000;
			{8'd26, 8'd24}: color_data = 12'h000;
			{8'd26, 8'd25}: color_data = 12'h000;
			{8'd26, 8'd26}: color_data = 12'h000;
			{8'd26, 8'd27}: color_data = 12'h000;
			{8'd26, 8'd28}: color_data = 12'h000;
			{8'd26, 8'd29}: color_data = 12'h000;
			{8'd26, 8'd30}: color_data = 12'h000;
			{8'd26, 8'd31}: color_data = 12'h000;
			{8'd26, 8'd32}: color_data = 12'h000;
			{8'd26, 8'd33}: color_data = 12'h610;
			{8'd26, 8'd34}: color_data = 12'he21;
			{8'd26, 8'd35}: color_data = 12'he21;
			{8'd26, 8'd36}: color_data = 12'he21;
			{8'd26, 8'd37}: color_data = 12'he21;
			{8'd26, 8'd38}: color_data = 12'he21;
			{8'd26, 8'd39}: color_data = 12'he21;
			{8'd26, 8'd40}: color_data = 12'he21;
			{8'd26, 8'd41}: color_data = 12'he21;
			{8'd26, 8'd42}: color_data = 12'he21;
			{8'd26, 8'd43}: color_data = 12'he21;
			{8'd26, 8'd44}: color_data = 12'he21;
			{8'd26, 8'd45}: color_data = 12'he21;
			{8'd26, 8'd46}: color_data = 12'he21;
			{8'd26, 8'd47}: color_data = 12'he21;
			{8'd26, 8'd48}: color_data = 12'he21;
			{8'd26, 8'd49}: color_data = 12'he21;
			{8'd26, 8'd50}: color_data = 12'ha10;
			{8'd26, 8'd51}: color_data = 12'h200;
			{8'd26, 8'd52}: color_data = 12'h000;
			{8'd26, 8'd53}: color_data = 12'h000;
			{8'd26, 8'd54}: color_data = 12'h000;
			{8'd26, 8'd55}: color_data = 12'h000;
			{8'd26, 8'd56}: color_data = 12'h000;
			{8'd26, 8'd57}: color_data = 12'h000;
			{8'd26, 8'd58}: color_data = 12'h000;
			{8'd26, 8'd59}: color_data = 12'h000;
			{8'd26, 8'd60}: color_data = 12'h000;
			{8'd26, 8'd61}: color_data = 12'h000;
			{8'd26, 8'd62}: color_data = 12'h000;
			{8'd26, 8'd63}: color_data = 12'h000;
			{8'd26, 8'd101}: color_data = 12'he00;
			{8'd26, 8'd102}: color_data = 12'he00;
			{8'd26, 8'd103}: color_data = 12'he00;
			{8'd26, 8'd104}: color_data = 12'he00;
			{8'd26, 8'd105}: color_data = 12'he00;
			{8'd26, 8'd106}: color_data = 12'he01;
			{8'd26, 8'd107}: color_data = 12'he00;
			{8'd26, 8'd136}: color_data = 12'he01;
			{8'd26, 8'd137}: color_data = 12'he00;
			{8'd26, 8'd138}: color_data = 12'he00;
			{8'd26, 8'd139}: color_data = 12'he00;
			{8'd26, 8'd140}: color_data = 12'he00;
			{8'd26, 8'd141}: color_data = 12'he00;
			{8'd26, 8'd142}: color_data = 12'he00;
			{8'd26, 8'd143}: color_data = 12'he01;
			{8'd27, 8'd8}: color_data = 12'h000;
			{8'd27, 8'd9}: color_data = 12'h000;
			{8'd27, 8'd10}: color_data = 12'h000;
			{8'd27, 8'd11}: color_data = 12'h000;
			{8'd27, 8'd12}: color_data = 12'h000;
			{8'd27, 8'd13}: color_data = 12'h000;
			{8'd27, 8'd14}: color_data = 12'h000;
			{8'd27, 8'd15}: color_data = 12'h000;
			{8'd27, 8'd16}: color_data = 12'h000;
			{8'd27, 8'd17}: color_data = 12'h000;
			{8'd27, 8'd19}: color_data = 12'h000;
			{8'd27, 8'd20}: color_data = 12'h000;
			{8'd27, 8'd21}: color_data = 12'h000;
			{8'd27, 8'd22}: color_data = 12'h001;
			{8'd27, 8'd23}: color_data = 12'h034;
			{8'd27, 8'd24}: color_data = 12'h000;
			{8'd27, 8'd25}: color_data = 12'h000;
			{8'd27, 8'd26}: color_data = 12'h000;
			{8'd27, 8'd27}: color_data = 12'h000;
			{8'd27, 8'd28}: color_data = 12'h000;
			{8'd27, 8'd29}: color_data = 12'h000;
			{8'd27, 8'd30}: color_data = 12'h000;
			{8'd27, 8'd31}: color_data = 12'h000;
			{8'd27, 8'd32}: color_data = 12'h000;
			{8'd27, 8'd33}: color_data = 12'h400;
			{8'd27, 8'd34}: color_data = 12'he21;
			{8'd27, 8'd35}: color_data = 12'he21;
			{8'd27, 8'd36}: color_data = 12'he21;
			{8'd27, 8'd37}: color_data = 12'he21;
			{8'd27, 8'd38}: color_data = 12'he21;
			{8'd27, 8'd39}: color_data = 12'he21;
			{8'd27, 8'd40}: color_data = 12'he21;
			{8'd27, 8'd41}: color_data = 12'he21;
			{8'd27, 8'd42}: color_data = 12'he21;
			{8'd27, 8'd43}: color_data = 12'he21;
			{8'd27, 8'd44}: color_data = 12'he21;
			{8'd27, 8'd45}: color_data = 12'he21;
			{8'd27, 8'd46}: color_data = 12'he21;
			{8'd27, 8'd47}: color_data = 12'he21;
			{8'd27, 8'd48}: color_data = 12'he21;
			{8'd27, 8'd49}: color_data = 12'he21;
			{8'd27, 8'd50}: color_data = 12'he21;
			{8'd27, 8'd51}: color_data = 12'hd20;
			{8'd27, 8'd52}: color_data = 12'h810;
			{8'd27, 8'd53}: color_data = 12'h100;
			{8'd27, 8'd54}: color_data = 12'h000;
			{8'd27, 8'd55}: color_data = 12'h000;
			{8'd27, 8'd56}: color_data = 12'h000;
			{8'd27, 8'd57}: color_data = 12'h000;
			{8'd27, 8'd58}: color_data = 12'h000;
			{8'd27, 8'd59}: color_data = 12'h000;
			{8'd27, 8'd60}: color_data = 12'h000;
			{8'd27, 8'd61}: color_data = 12'h000;
			{8'd27, 8'd62}: color_data = 12'h000;
			{8'd27, 8'd63}: color_data = 12'h000;
			{8'd27, 8'd101}: color_data = 12'he00;
			{8'd27, 8'd102}: color_data = 12'he01;
			{8'd27, 8'd103}: color_data = 12'he00;
			{8'd27, 8'd104}: color_data = 12'he00;
			{8'd27, 8'd105}: color_data = 12'he00;
			{8'd27, 8'd106}: color_data = 12'he00;
			{8'd27, 8'd107}: color_data = 12'he00;
			{8'd27, 8'd137}: color_data = 12'he00;
			{8'd27, 8'd138}: color_data = 12'he00;
			{8'd27, 8'd139}: color_data = 12'he00;
			{8'd27, 8'd140}: color_data = 12'he00;
			{8'd27, 8'd141}: color_data = 12'he00;
			{8'd27, 8'd142}: color_data = 12'he00;
			{8'd27, 8'd143}: color_data = 12'he00;
			{8'd28, 8'd7}: color_data = 12'h000;
			{8'd28, 8'd8}: color_data = 12'h000;
			{8'd28, 8'd9}: color_data = 12'h000;
			{8'd28, 8'd10}: color_data = 12'h000;
			{8'd28, 8'd11}: color_data = 12'h023;
			{8'd28, 8'd12}: color_data = 12'h001;
			{8'd28, 8'd13}: color_data = 12'h000;
			{8'd28, 8'd14}: color_data = 12'h000;
			{8'd28, 8'd15}: color_data = 12'h000;
			{8'd28, 8'd16}: color_data = 12'h000;
			{8'd28, 8'd17}: color_data = 12'h000;
			{8'd28, 8'd18}: color_data = 12'h000;
			{8'd28, 8'd19}: color_data = 12'h000;
			{8'd28, 8'd20}: color_data = 12'h000;
			{8'd28, 8'd21}: color_data = 12'h012;
			{8'd28, 8'd22}: color_data = 12'h07a;
			{8'd28, 8'd23}: color_data = 12'h0ae;
			{8'd28, 8'd24}: color_data = 12'h046;
			{8'd28, 8'd25}: color_data = 12'h000;
			{8'd28, 8'd26}: color_data = 12'h000;
			{8'd28, 8'd27}: color_data = 12'h000;
			{8'd28, 8'd28}: color_data = 12'h000;
			{8'd28, 8'd29}: color_data = 12'h000;
			{8'd28, 8'd30}: color_data = 12'h000;
			{8'd28, 8'd31}: color_data = 12'h000;
			{8'd28, 8'd32}: color_data = 12'h000;
			{8'd28, 8'd33}: color_data = 12'h200;
			{8'd28, 8'd34}: color_data = 12'he21;
			{8'd28, 8'd35}: color_data = 12'he21;
			{8'd28, 8'd36}: color_data = 12'he21;
			{8'd28, 8'd37}: color_data = 12'he21;
			{8'd28, 8'd38}: color_data = 12'he21;
			{8'd28, 8'd39}: color_data = 12'he21;
			{8'd28, 8'd40}: color_data = 12'he21;
			{8'd28, 8'd41}: color_data = 12'he21;
			{8'd28, 8'd42}: color_data = 12'he21;
			{8'd28, 8'd43}: color_data = 12'he21;
			{8'd28, 8'd44}: color_data = 12'he21;
			{8'd28, 8'd45}: color_data = 12'he21;
			{8'd28, 8'd46}: color_data = 12'he21;
			{8'd28, 8'd47}: color_data = 12'he21;
			{8'd28, 8'd48}: color_data = 12'he21;
			{8'd28, 8'd49}: color_data = 12'he21;
			{8'd28, 8'd50}: color_data = 12'he21;
			{8'd28, 8'd51}: color_data = 12'he21;
			{8'd28, 8'd52}: color_data = 12'he21;
			{8'd28, 8'd53}: color_data = 12'hd20;
			{8'd28, 8'd54}: color_data = 12'h610;
			{8'd28, 8'd55}: color_data = 12'h000;
			{8'd28, 8'd56}: color_data = 12'h000;
			{8'd28, 8'd57}: color_data = 12'h000;
			{8'd28, 8'd58}: color_data = 12'h000;
			{8'd28, 8'd59}: color_data = 12'h000;
			{8'd28, 8'd60}: color_data = 12'h000;
			{8'd28, 8'd61}: color_data = 12'h000;
			{8'd28, 8'd62}: color_data = 12'h000;
			{8'd28, 8'd63}: color_data = 12'h000;
			{8'd28, 8'd64}: color_data = 12'h000;
			{8'd28, 8'd100}: color_data = 12'hf00;
			{8'd28, 8'd101}: color_data = 12'he00;
			{8'd28, 8'd102}: color_data = 12'he00;
			{8'd28, 8'd103}: color_data = 12'he00;
			{8'd28, 8'd104}: color_data = 12'he00;
			{8'd28, 8'd105}: color_data = 12'he00;
			{8'd28, 8'd106}: color_data = 12'he00;
			{8'd28, 8'd107}: color_data = 12'hd00;
			{8'd28, 8'd137}: color_data = 12'he00;
			{8'd28, 8'd138}: color_data = 12'he00;
			{8'd28, 8'd139}: color_data = 12'he00;
			{8'd28, 8'd140}: color_data = 12'he00;
			{8'd28, 8'd141}: color_data = 12'he00;
			{8'd28, 8'd142}: color_data = 12'he01;
			{8'd28, 8'd143}: color_data = 12'he00;
			{8'd29, 8'd5}: color_data = 12'h000;
			{8'd29, 8'd6}: color_data = 12'h000;
			{8'd29, 8'd7}: color_data = 12'h000;
			{8'd29, 8'd8}: color_data = 12'h000;
			{8'd29, 8'd9}: color_data = 12'h001;
			{8'd29, 8'd10}: color_data = 12'h058;
			{8'd29, 8'd11}: color_data = 12'h0ae;
			{8'd29, 8'd12}: color_data = 12'h057;
			{8'd29, 8'd13}: color_data = 12'h000;
			{8'd29, 8'd14}: color_data = 12'h000;
			{8'd29, 8'd15}: color_data = 12'h000;
			{8'd29, 8'd16}: color_data = 12'h000;
			{8'd29, 8'd17}: color_data = 12'h000;
			{8'd29, 8'd18}: color_data = 12'h000;
			{8'd29, 8'd19}: color_data = 12'h000;
			{8'd29, 8'd20}: color_data = 12'h034;
			{8'd29, 8'd21}: color_data = 12'h09c;
			{8'd29, 8'd22}: color_data = 12'h0ae;
			{8'd29, 8'd23}: color_data = 12'h09d;
			{8'd29, 8'd24}: color_data = 12'h09d;
			{8'd29, 8'd25}: color_data = 12'h035;
			{8'd29, 8'd26}: color_data = 12'h000;
			{8'd29, 8'd27}: color_data = 12'h000;
			{8'd29, 8'd28}: color_data = 12'h000;
			{8'd29, 8'd29}: color_data = 12'h000;
			{8'd29, 8'd30}: color_data = 12'h000;
			{8'd29, 8'd31}: color_data = 12'h000;
			{8'd29, 8'd32}: color_data = 12'h000;
			{8'd29, 8'd33}: color_data = 12'h000;
			{8'd29, 8'd34}: color_data = 12'h500;
			{8'd29, 8'd35}: color_data = 12'ha10;
			{8'd29, 8'd36}: color_data = 12'hd20;
			{8'd29, 8'd37}: color_data = 12'he21;
			{8'd29, 8'd38}: color_data = 12'he21;
			{8'd29, 8'd39}: color_data = 12'he21;
			{8'd29, 8'd40}: color_data = 12'he21;
			{8'd29, 8'd41}: color_data = 12'he21;
			{8'd29, 8'd42}: color_data = 12'he21;
			{8'd29, 8'd43}: color_data = 12'he21;
			{8'd29, 8'd44}: color_data = 12'he21;
			{8'd29, 8'd45}: color_data = 12'he21;
			{8'd29, 8'd46}: color_data = 12'he21;
			{8'd29, 8'd47}: color_data = 12'he21;
			{8'd29, 8'd48}: color_data = 12'he21;
			{8'd29, 8'd49}: color_data = 12'he21;
			{8'd29, 8'd50}: color_data = 12'he21;
			{8'd29, 8'd51}: color_data = 12'he21;
			{8'd29, 8'd52}: color_data = 12'he21;
			{8'd29, 8'd53}: color_data = 12'he21;
			{8'd29, 8'd54}: color_data = 12'he21;
			{8'd29, 8'd55}: color_data = 12'hc10;
			{8'd29, 8'd56}: color_data = 12'h500;
			{8'd29, 8'd57}: color_data = 12'h000;
			{8'd29, 8'd58}: color_data = 12'h000;
			{8'd29, 8'd59}: color_data = 12'h000;
			{8'd29, 8'd60}: color_data = 12'h000;
			{8'd29, 8'd61}: color_data = 12'h000;
			{8'd29, 8'd62}: color_data = 12'h000;
			{8'd29, 8'd63}: color_data = 12'h000;
			{8'd29, 8'd64}: color_data = 12'h000;
			{8'd29, 8'd65}: color_data = 12'h000;
			{8'd29, 8'd66}: color_data = 12'h000;
			{8'd29, 8'd100}: color_data = 12'he00;
			{8'd29, 8'd101}: color_data = 12'he00;
			{8'd29, 8'd102}: color_data = 12'he00;
			{8'd29, 8'd103}: color_data = 12'he00;
			{8'd29, 8'd104}: color_data = 12'he00;
			{8'd29, 8'd105}: color_data = 12'he01;
			{8'd29, 8'd106}: color_data = 12'he00;
			{8'd29, 8'd111}: color_data = 12'hd00;
			{8'd29, 8'd112}: color_data = 12'he00;
			{8'd29, 8'd113}: color_data = 12'hf00;
			{8'd29, 8'd138}: color_data = 12'he00;
			{8'd29, 8'd139}: color_data = 12'he01;
			{8'd29, 8'd140}: color_data = 12'he00;
			{8'd29, 8'd141}: color_data = 12'he00;
			{8'd29, 8'd142}: color_data = 12'he00;
			{8'd29, 8'd143}: color_data = 12'he00;
			{8'd29, 8'd144}: color_data = 12'he01;
			{8'd30, 8'd4}: color_data = 12'h000;
			{8'd30, 8'd5}: color_data = 12'h000;
			{8'd30, 8'd6}: color_data = 12'h000;
			{8'd30, 8'd7}: color_data = 12'h000;
			{8'd30, 8'd8}: color_data = 12'h024;
			{8'd30, 8'd9}: color_data = 12'h08b;
			{8'd30, 8'd10}: color_data = 12'h0ae;
			{8'd30, 8'd11}: color_data = 12'h09d;
			{8'd30, 8'd12}: color_data = 12'h09d;
			{8'd30, 8'd13}: color_data = 12'h012;
			{8'd30, 8'd14}: color_data = 12'h000;
			{8'd30, 8'd15}: color_data = 12'h000;
			{8'd30, 8'd16}: color_data = 12'h000;
			{8'd30, 8'd17}: color_data = 12'h000;
			{8'd30, 8'd18}: color_data = 12'h000;
			{8'd30, 8'd19}: color_data = 12'h057;
			{8'd30, 8'd20}: color_data = 12'h09d;
			{8'd30, 8'd21}: color_data = 12'h09d;
			{8'd30, 8'd22}: color_data = 12'h09d;
			{8'd30, 8'd23}: color_data = 12'h09d;
			{8'd30, 8'd24}: color_data = 12'h09d;
			{8'd30, 8'd25}: color_data = 12'h09d;
			{8'd30, 8'd26}: color_data = 12'h023;
			{8'd30, 8'd27}: color_data = 12'h000;
			{8'd30, 8'd28}: color_data = 12'h000;
			{8'd30, 8'd29}: color_data = 12'h000;
			{8'd30, 8'd30}: color_data = 12'h000;
			{8'd30, 8'd31}: color_data = 12'h000;
			{8'd30, 8'd32}: color_data = 12'h000;
			{8'd30, 8'd33}: color_data = 12'h000;
			{8'd30, 8'd34}: color_data = 12'h000;
			{8'd30, 8'd35}: color_data = 12'h000;
			{8'd30, 8'd36}: color_data = 12'h100;
			{8'd30, 8'd37}: color_data = 12'h500;
			{8'd30, 8'd38}: color_data = 12'ha10;
			{8'd30, 8'd39}: color_data = 12'hd20;
			{8'd30, 8'd40}: color_data = 12'he21;
			{8'd30, 8'd41}: color_data = 12'he21;
			{8'd30, 8'd42}: color_data = 12'he21;
			{8'd30, 8'd43}: color_data = 12'he21;
			{8'd30, 8'd44}: color_data = 12'he21;
			{8'd30, 8'd45}: color_data = 12'he21;
			{8'd30, 8'd46}: color_data = 12'he21;
			{8'd30, 8'd47}: color_data = 12'he21;
			{8'd30, 8'd48}: color_data = 12'he21;
			{8'd30, 8'd49}: color_data = 12'he21;
			{8'd30, 8'd50}: color_data = 12'he21;
			{8'd30, 8'd51}: color_data = 12'he21;
			{8'd30, 8'd52}: color_data = 12'he21;
			{8'd30, 8'd53}: color_data = 12'he21;
			{8'd30, 8'd54}: color_data = 12'he21;
			{8'd30, 8'd55}: color_data = 12'he21;
			{8'd30, 8'd56}: color_data = 12'he21;
			{8'd30, 8'd57}: color_data = 12'ha10;
			{8'd30, 8'd58}: color_data = 12'h300;
			{8'd30, 8'd59}: color_data = 12'h000;
			{8'd30, 8'd60}: color_data = 12'h000;
			{8'd30, 8'd61}: color_data = 12'h000;
			{8'd30, 8'd62}: color_data = 12'h000;
			{8'd30, 8'd63}: color_data = 12'h000;
			{8'd30, 8'd64}: color_data = 12'h000;
			{8'd30, 8'd65}: color_data = 12'h000;
			{8'd30, 8'd66}: color_data = 12'h000;
			{8'd30, 8'd67}: color_data = 12'h000;
			{8'd30, 8'd68}: color_data = 12'h000;
			{8'd30, 8'd100}: color_data = 12'he00;
			{8'd30, 8'd101}: color_data = 12'he00;
			{8'd30, 8'd102}: color_data = 12'he00;
			{8'd30, 8'd103}: color_data = 12'he00;
			{8'd30, 8'd104}: color_data = 12'he00;
			{8'd30, 8'd105}: color_data = 12'he00;
			{8'd30, 8'd106}: color_data = 12'he00;
			{8'd30, 8'd111}: color_data = 12'he00;
			{8'd30, 8'd112}: color_data = 12'he00;
			{8'd30, 8'd113}: color_data = 12'he00;
			{8'd30, 8'd114}: color_data = 12'he00;
			{8'd30, 8'd115}: color_data = 12'he00;
			{8'd30, 8'd138}: color_data = 12'he00;
			{8'd30, 8'd139}: color_data = 12'he01;
			{8'd30, 8'd140}: color_data = 12'he00;
			{8'd30, 8'd141}: color_data = 12'he00;
			{8'd30, 8'd142}: color_data = 12'he00;
			{8'd30, 8'd143}: color_data = 12'he00;
			{8'd30, 8'd144}: color_data = 12'he00;
			{8'd31, 8'd2}: color_data = 12'h000;
			{8'd31, 8'd3}: color_data = 12'h000;
			{8'd31, 8'd4}: color_data = 12'h000;
			{8'd31, 8'd5}: color_data = 12'h000;
			{8'd31, 8'd6}: color_data = 12'h001;
			{8'd31, 8'd7}: color_data = 12'h058;
			{8'd31, 8'd8}: color_data = 12'h09d;
			{8'd31, 8'd9}: color_data = 12'h09d;
			{8'd31, 8'd10}: color_data = 12'h09d;
			{8'd31, 8'd11}: color_data = 12'h09d;
			{8'd31, 8'd12}: color_data = 12'h0ae;
			{8'd31, 8'd13}: color_data = 12'h079;
			{8'd31, 8'd14}: color_data = 12'h000;
			{8'd31, 8'd15}: color_data = 12'h000;
			{8'd31, 8'd16}: color_data = 12'h000;
			{8'd31, 8'd17}: color_data = 12'h011;
			{8'd31, 8'd18}: color_data = 12'h07a;
			{8'd31, 8'd19}: color_data = 12'h0ae;
			{8'd31, 8'd20}: color_data = 12'h09d;
			{8'd31, 8'd21}: color_data = 12'h09d;
			{8'd31, 8'd22}: color_data = 12'h09d;
			{8'd31, 8'd23}: color_data = 12'h09d;
			{8'd31, 8'd24}: color_data = 12'h09d;
			{8'd31, 8'd25}: color_data = 12'h09d;
			{8'd31, 8'd26}: color_data = 12'h08c;
			{8'd31, 8'd27}: color_data = 12'h012;
			{8'd31, 8'd28}: color_data = 12'h000;
			{8'd31, 8'd29}: color_data = 12'h000;
			{8'd31, 8'd30}: color_data = 12'h000;
			{8'd31, 8'd31}: color_data = 12'h000;
			{8'd31, 8'd32}: color_data = 12'h000;
			{8'd31, 8'd33}: color_data = 12'h000;
			{8'd31, 8'd34}: color_data = 12'h000;
			{8'd31, 8'd35}: color_data = 12'h000;
			{8'd31, 8'd36}: color_data = 12'h000;
			{8'd31, 8'd37}: color_data = 12'h000;
			{8'd31, 8'd38}: color_data = 12'h000;
			{8'd31, 8'd39}: color_data = 12'h100;
			{8'd31, 8'd40}: color_data = 12'h500;
			{8'd31, 8'd41}: color_data = 12'ha10;
			{8'd31, 8'd42}: color_data = 12'hd20;
			{8'd31, 8'd43}: color_data = 12'he21;
			{8'd31, 8'd44}: color_data = 12'he21;
			{8'd31, 8'd45}: color_data = 12'he21;
			{8'd31, 8'd46}: color_data = 12'he21;
			{8'd31, 8'd47}: color_data = 12'he21;
			{8'd31, 8'd48}: color_data = 12'he21;
			{8'd31, 8'd49}: color_data = 12'he21;
			{8'd31, 8'd50}: color_data = 12'he21;
			{8'd31, 8'd51}: color_data = 12'he21;
			{8'd31, 8'd52}: color_data = 12'he21;
			{8'd31, 8'd53}: color_data = 12'he21;
			{8'd31, 8'd54}: color_data = 12'he21;
			{8'd31, 8'd55}: color_data = 12'he21;
			{8'd31, 8'd56}: color_data = 12'he21;
			{8'd31, 8'd57}: color_data = 12'hf21;
			{8'd31, 8'd58}: color_data = 12'hd20;
			{8'd31, 8'd59}: color_data = 12'h100;
			{8'd31, 8'd60}: color_data = 12'h000;
			{8'd31, 8'd61}: color_data = 12'h000;
			{8'd31, 8'd62}: color_data = 12'h000;
			{8'd31, 8'd63}: color_data = 12'h000;
			{8'd31, 8'd64}: color_data = 12'h000;
			{8'd31, 8'd65}: color_data = 12'h000;
			{8'd31, 8'd66}: color_data = 12'h000;
			{8'd31, 8'd67}: color_data = 12'h000;
			{8'd31, 8'd68}: color_data = 12'h000;
			{8'd31, 8'd100}: color_data = 12'he00;
			{8'd31, 8'd101}: color_data = 12'he01;
			{8'd31, 8'd102}: color_data = 12'he00;
			{8'd31, 8'd103}: color_data = 12'he00;
			{8'd31, 8'd104}: color_data = 12'he00;
			{8'd31, 8'd105}: color_data = 12'he00;
			{8'd31, 8'd106}: color_data = 12'he00;
			{8'd31, 8'd111}: color_data = 12'he00;
			{8'd31, 8'd112}: color_data = 12'he00;
			{8'd31, 8'd113}: color_data = 12'he00;
			{8'd31, 8'd114}: color_data = 12'he01;
			{8'd31, 8'd115}: color_data = 12'he00;
			{8'd31, 8'd116}: color_data = 12'he00;
			{8'd31, 8'd117}: color_data = 12'he01;
			{8'd31, 8'd118}: color_data = 12'he00;
			{8'd31, 8'd138}: color_data = 12'he00;
			{8'd31, 8'd139}: color_data = 12'he00;
			{8'd31, 8'd140}: color_data = 12'he00;
			{8'd31, 8'd141}: color_data = 12'he00;
			{8'd31, 8'd142}: color_data = 12'he00;
			{8'd31, 8'd143}: color_data = 12'he00;
			{8'd31, 8'd144}: color_data = 12'he00;
			{8'd32, 8'd1}: color_data = 12'h000;
			{8'd32, 8'd2}: color_data = 12'h000;
			{8'd32, 8'd3}: color_data = 12'h000;
			{8'd32, 8'd4}: color_data = 12'h000;
			{8'd32, 8'd5}: color_data = 12'h023;
			{8'd32, 8'd6}: color_data = 12'h08b;
			{8'd32, 8'd7}: color_data = 12'h0ae;
			{8'd32, 8'd8}: color_data = 12'h09d;
			{8'd32, 8'd9}: color_data = 12'h09d;
			{8'd32, 8'd10}: color_data = 12'h09d;
			{8'd32, 8'd11}: color_data = 12'h09d;
			{8'd32, 8'd12}: color_data = 12'h09d;
			{8'd32, 8'd13}: color_data = 12'h09d;
			{8'd32, 8'd14}: color_data = 12'h035;
			{8'd32, 8'd15}: color_data = 12'h000;
			{8'd32, 8'd16}: color_data = 12'h000;
			{8'd32, 8'd17}: color_data = 12'h011;
			{8'd32, 8'd18}: color_data = 12'h08b;
			{8'd32, 8'd19}: color_data = 12'h09d;
			{8'd32, 8'd20}: color_data = 12'h09d;
			{8'd32, 8'd21}: color_data = 12'h09d;
			{8'd32, 8'd22}: color_data = 12'h09d;
			{8'd32, 8'd23}: color_data = 12'h09d;
			{8'd32, 8'd24}: color_data = 12'h09d;
			{8'd32, 8'd25}: color_data = 12'h09d;
			{8'd32, 8'd26}: color_data = 12'h0ae;
			{8'd32, 8'd27}: color_data = 12'h07b;
			{8'd32, 8'd28}: color_data = 12'h001;
			{8'd32, 8'd29}: color_data = 12'h000;
			{8'd32, 8'd30}: color_data = 12'h000;
			{8'd32, 8'd31}: color_data = 12'h000;
			{8'd32, 8'd32}: color_data = 12'h000;
			{8'd32, 8'd33}: color_data = 12'h000;
			{8'd32, 8'd34}: color_data = 12'h000;
			{8'd32, 8'd35}: color_data = 12'h000;
			{8'd32, 8'd36}: color_data = 12'h000;
			{8'd32, 8'd37}: color_data = 12'h000;
			{8'd32, 8'd38}: color_data = 12'h000;
			{8'd32, 8'd39}: color_data = 12'h000;
			{8'd32, 8'd40}: color_data = 12'h000;
			{8'd32, 8'd41}: color_data = 12'h000;
			{8'd32, 8'd42}: color_data = 12'h100;
			{8'd32, 8'd43}: color_data = 12'h500;
			{8'd32, 8'd44}: color_data = 12'hc10;
			{8'd32, 8'd45}: color_data = 12'he21;
			{8'd32, 8'd46}: color_data = 12'he21;
			{8'd32, 8'd47}: color_data = 12'he21;
			{8'd32, 8'd48}: color_data = 12'he21;
			{8'd32, 8'd49}: color_data = 12'he21;
			{8'd32, 8'd50}: color_data = 12'he21;
			{8'd32, 8'd51}: color_data = 12'he21;
			{8'd32, 8'd52}: color_data = 12'he21;
			{8'd32, 8'd53}: color_data = 12'he21;
			{8'd32, 8'd54}: color_data = 12'he21;
			{8'd32, 8'd55}: color_data = 12'he21;
			{8'd32, 8'd56}: color_data = 12'he21;
			{8'd32, 8'd57}: color_data = 12'hc10;
			{8'd32, 8'd58}: color_data = 12'h300;
			{8'd32, 8'd59}: color_data = 12'h000;
			{8'd32, 8'd60}: color_data = 12'h000;
			{8'd32, 8'd61}: color_data = 12'h000;
			{8'd32, 8'd62}: color_data = 12'h000;
			{8'd32, 8'd63}: color_data = 12'h000;
			{8'd32, 8'd64}: color_data = 12'h000;
			{8'd32, 8'd65}: color_data = 12'h000;
			{8'd32, 8'd66}: color_data = 12'h000;
			{8'd32, 8'd100}: color_data = 12'he00;
			{8'd32, 8'd101}: color_data = 12'he01;
			{8'd32, 8'd102}: color_data = 12'he00;
			{8'd32, 8'd103}: color_data = 12'he00;
			{8'd32, 8'd104}: color_data = 12'he00;
			{8'd32, 8'd105}: color_data = 12'he00;
			{8'd32, 8'd106}: color_data = 12'he00;
			{8'd32, 8'd111}: color_data = 12'he01;
			{8'd32, 8'd112}: color_data = 12'he00;
			{8'd32, 8'd113}: color_data = 12'he00;
			{8'd32, 8'd114}: color_data = 12'he00;
			{8'd32, 8'd115}: color_data = 12'he00;
			{8'd32, 8'd116}: color_data = 12'he01;
			{8'd32, 8'd117}: color_data = 12'he01;
			{8'd32, 8'd118}: color_data = 12'he00;
			{8'd32, 8'd119}: color_data = 12'he00;
			{8'd32, 8'd120}: color_data = 12'he01;
			{8'd32, 8'd121}: color_data = 12'hd00;
			{8'd32, 8'd138}: color_data = 12'he00;
			{8'd32, 8'd139}: color_data = 12'he00;
			{8'd32, 8'd140}: color_data = 12'he00;
			{8'd32, 8'd141}: color_data = 12'he00;
			{8'd32, 8'd142}: color_data = 12'he00;
			{8'd32, 8'd143}: color_data = 12'he00;
			{8'd32, 8'd144}: color_data = 12'he00;
			{8'd33, 8'd0}: color_data = 12'h000;
			{8'd33, 8'd1}: color_data = 12'h000;
			{8'd33, 8'd2}: color_data = 12'h000;
			{8'd33, 8'd3}: color_data = 12'h000;
			{8'd33, 8'd4}: color_data = 12'h057;
			{8'd33, 8'd5}: color_data = 12'h09d;
			{8'd33, 8'd6}: color_data = 12'h09d;
			{8'd33, 8'd7}: color_data = 12'h09d;
			{8'd33, 8'd8}: color_data = 12'h09d;
			{8'd33, 8'd9}: color_data = 12'h09d;
			{8'd33, 8'd10}: color_data = 12'h09d;
			{8'd33, 8'd11}: color_data = 12'h09d;
			{8'd33, 8'd12}: color_data = 12'h09d;
			{8'd33, 8'd13}: color_data = 12'h09d;
			{8'd33, 8'd14}: color_data = 12'h08c;
			{8'd33, 8'd15}: color_data = 12'h001;
			{8'd33, 8'd16}: color_data = 12'h000;
			{8'd33, 8'd17}: color_data = 12'h000;
			{8'd33, 8'd18}: color_data = 12'h022;
			{8'd33, 8'd19}: color_data = 12'h09c;
			{8'd33, 8'd20}: color_data = 12'h09d;
			{8'd33, 8'd21}: color_data = 12'h09d;
			{8'd33, 8'd22}: color_data = 12'h09d;
			{8'd33, 8'd23}: color_data = 12'h09d;
			{8'd33, 8'd24}: color_data = 12'h09d;
			{8'd33, 8'd25}: color_data = 12'h09d;
			{8'd33, 8'd26}: color_data = 12'h09d;
			{8'd33, 8'd27}: color_data = 12'h0ae;
			{8'd33, 8'd28}: color_data = 12'h069;
			{8'd33, 8'd29}: color_data = 12'h000;
			{8'd33, 8'd30}: color_data = 12'h000;
			{8'd33, 8'd31}: color_data = 12'h000;
			{8'd33, 8'd32}: color_data = 12'h000;
			{8'd33, 8'd33}: color_data = 12'h000;
			{8'd33, 8'd34}: color_data = 12'h000;
			{8'd33, 8'd35}: color_data = 12'h000;
			{8'd33, 8'd36}: color_data = 12'h000;
			{8'd33, 8'd37}: color_data = 12'h000;
			{8'd33, 8'd38}: color_data = 12'h000;
			{8'd33, 8'd39}: color_data = 12'h000;
			{8'd33, 8'd40}: color_data = 12'h000;
			{8'd33, 8'd41}: color_data = 12'h000;
			{8'd33, 8'd42}: color_data = 12'h100;
			{8'd33, 8'd43}: color_data = 12'h710;
			{8'd33, 8'd44}: color_data = 12'hd20;
			{8'd33, 8'd45}: color_data = 12'he21;
			{8'd33, 8'd46}: color_data = 12'he21;
			{8'd33, 8'd47}: color_data = 12'he21;
			{8'd33, 8'd48}: color_data = 12'he21;
			{8'd33, 8'd49}: color_data = 12'he21;
			{8'd33, 8'd50}: color_data = 12'he21;
			{8'd33, 8'd51}: color_data = 12'he21;
			{8'd33, 8'd52}: color_data = 12'he21;
			{8'd33, 8'd53}: color_data = 12'he21;
			{8'd33, 8'd54}: color_data = 12'he21;
			{8'd33, 8'd55}: color_data = 12'he21;
			{8'd33, 8'd56}: color_data = 12'ha10;
			{8'd33, 8'd57}: color_data = 12'h100;
			{8'd33, 8'd58}: color_data = 12'h000;
			{8'd33, 8'd59}: color_data = 12'h000;
			{8'd33, 8'd60}: color_data = 12'h000;
			{8'd33, 8'd61}: color_data = 12'h000;
			{8'd33, 8'd62}: color_data = 12'h000;
			{8'd33, 8'd63}: color_data = 12'h000;
			{8'd33, 8'd64}: color_data = 12'h000;
			{8'd33, 8'd65}: color_data = 12'h000;
			{8'd33, 8'd100}: color_data = 12'he00;
			{8'd33, 8'd101}: color_data = 12'he01;
			{8'd33, 8'd102}: color_data = 12'he00;
			{8'd33, 8'd103}: color_data = 12'he00;
			{8'd33, 8'd104}: color_data = 12'he00;
			{8'd33, 8'd105}: color_data = 12'he00;
			{8'd33, 8'd106}: color_data = 12'he01;
			{8'd33, 8'd111}: color_data = 12'he01;
			{8'd33, 8'd112}: color_data = 12'he00;
			{8'd33, 8'd113}: color_data = 12'he00;
			{8'd33, 8'd114}: color_data = 12'he00;
			{8'd33, 8'd115}: color_data = 12'he00;
			{8'd33, 8'd116}: color_data = 12'he00;
			{8'd33, 8'd117}: color_data = 12'he00;
			{8'd33, 8'd118}: color_data = 12'he00;
			{8'd33, 8'd119}: color_data = 12'he01;
			{8'd33, 8'd120}: color_data = 12'he00;
			{8'd33, 8'd121}: color_data = 12'he00;
			{8'd33, 8'd122}: color_data = 12'he00;
			{8'd33, 8'd123}: color_data = 12'he00;
			{8'd33, 8'd138}: color_data = 12'he01;
			{8'd33, 8'd139}: color_data = 12'he00;
			{8'd33, 8'd140}: color_data = 12'he00;
			{8'd33, 8'd141}: color_data = 12'he00;
			{8'd33, 8'd142}: color_data = 12'he00;
			{8'd33, 8'd143}: color_data = 12'he01;
			{8'd33, 8'd144}: color_data = 12'he00;
			{8'd34, 8'd0}: color_data = 12'h000;
			{8'd34, 8'd1}: color_data = 12'h000;
			{8'd34, 8'd2}: color_data = 12'h000;
			{8'd34, 8'd3}: color_data = 12'h068;
			{8'd34, 8'd4}: color_data = 12'h0ae;
			{8'd34, 8'd5}: color_data = 12'h09d;
			{8'd34, 8'd6}: color_data = 12'h09d;
			{8'd34, 8'd7}: color_data = 12'h09d;
			{8'd34, 8'd8}: color_data = 12'h09d;
			{8'd34, 8'd9}: color_data = 12'h09d;
			{8'd34, 8'd10}: color_data = 12'h09d;
			{8'd34, 8'd11}: color_data = 12'h09d;
			{8'd34, 8'd12}: color_data = 12'h09d;
			{8'd34, 8'd13}: color_data = 12'h09d;
			{8'd34, 8'd14}: color_data = 12'h0ae;
			{8'd34, 8'd15}: color_data = 12'h057;
			{8'd34, 8'd16}: color_data = 12'h000;
			{8'd34, 8'd17}: color_data = 12'h000;
			{8'd34, 8'd18}: color_data = 12'h000;
			{8'd34, 8'd19}: color_data = 12'h034;
			{8'd34, 8'd20}: color_data = 12'h09d;
			{8'd34, 8'd21}: color_data = 12'h09d;
			{8'd34, 8'd22}: color_data = 12'h09d;
			{8'd34, 8'd23}: color_data = 12'h09d;
			{8'd34, 8'd24}: color_data = 12'h09d;
			{8'd34, 8'd25}: color_data = 12'h09d;
			{8'd34, 8'd26}: color_data = 12'h09d;
			{8'd34, 8'd27}: color_data = 12'h09d;
			{8'd34, 8'd28}: color_data = 12'h0ae;
			{8'd34, 8'd29}: color_data = 12'h058;
			{8'd34, 8'd30}: color_data = 12'h000;
			{8'd34, 8'd31}: color_data = 12'h000;
			{8'd34, 8'd32}: color_data = 12'h000;
			{8'd34, 8'd33}: color_data = 12'h000;
			{8'd34, 8'd34}: color_data = 12'h000;
			{8'd34, 8'd35}: color_data = 12'h000;
			{8'd34, 8'd36}: color_data = 12'h000;
			{8'd34, 8'd37}: color_data = 12'h000;
			{8'd34, 8'd38}: color_data = 12'h000;
			{8'd34, 8'd39}: color_data = 12'h000;
			{8'd34, 8'd40}: color_data = 12'h100;
			{8'd34, 8'd41}: color_data = 12'h710;
			{8'd34, 8'd42}: color_data = 12'hd20;
			{8'd34, 8'd43}: color_data = 12'he21;
			{8'd34, 8'd44}: color_data = 12'he21;
			{8'd34, 8'd45}: color_data = 12'he21;
			{8'd34, 8'd46}: color_data = 12'he21;
			{8'd34, 8'd47}: color_data = 12'he21;
			{8'd34, 8'd48}: color_data = 12'he21;
			{8'd34, 8'd49}: color_data = 12'he21;
			{8'd34, 8'd50}: color_data = 12'he21;
			{8'd34, 8'd51}: color_data = 12'he21;
			{8'd34, 8'd52}: color_data = 12'he21;
			{8'd34, 8'd53}: color_data = 12'he21;
			{8'd34, 8'd54}: color_data = 12'he21;
			{8'd34, 8'd55}: color_data = 12'h810;
			{8'd34, 8'd56}: color_data = 12'h000;
			{8'd34, 8'd57}: color_data = 12'h000;
			{8'd34, 8'd58}: color_data = 12'h000;
			{8'd34, 8'd59}: color_data = 12'h000;
			{8'd34, 8'd60}: color_data = 12'h000;
			{8'd34, 8'd61}: color_data = 12'h000;
			{8'd34, 8'd62}: color_data = 12'h000;
			{8'd34, 8'd63}: color_data = 12'h000;
			{8'd34, 8'd64}: color_data = 12'h000;
			{8'd34, 8'd100}: color_data = 12'he00;
			{8'd34, 8'd101}: color_data = 12'hf01;
			{8'd34, 8'd102}: color_data = 12'he00;
			{8'd34, 8'd103}: color_data = 12'he00;
			{8'd34, 8'd104}: color_data = 12'he00;
			{8'd34, 8'd105}: color_data = 12'he00;
			{8'd34, 8'd106}: color_data = 12'hc00;
			{8'd34, 8'd111}: color_data = 12'he01;
			{8'd34, 8'd112}: color_data = 12'he00;
			{8'd34, 8'd113}: color_data = 12'he00;
			{8'd34, 8'd114}: color_data = 12'he00;
			{8'd34, 8'd115}: color_data = 12'he00;
			{8'd34, 8'd116}: color_data = 12'he00;
			{8'd34, 8'd117}: color_data = 12'he00;
			{8'd34, 8'd118}: color_data = 12'he00;
			{8'd34, 8'd119}: color_data = 12'he00;
			{8'd34, 8'd120}: color_data = 12'he00;
			{8'd34, 8'd121}: color_data = 12'he00;
			{8'd34, 8'd122}: color_data = 12'he01;
			{8'd34, 8'd123}: color_data = 12'he00;
			{8'd34, 8'd124}: color_data = 12'he00;
			{8'd34, 8'd125}: color_data = 12'he00;
			{8'd34, 8'd126}: color_data = 12'hd00;
			{8'd34, 8'd138}: color_data = 12'he00;
			{8'd34, 8'd139}: color_data = 12'he00;
			{8'd34, 8'd140}: color_data = 12'he00;
			{8'd34, 8'd141}: color_data = 12'he00;
			{8'd34, 8'd142}: color_data = 12'he00;
			{8'd34, 8'd143}: color_data = 12'he01;
			{8'd34, 8'd144}: color_data = 12'he00;
			{8'd35, 8'd0}: color_data = 12'h000;
			{8'd35, 8'd1}: color_data = 12'h000;
			{8'd35, 8'd2}: color_data = 12'h000;
			{8'd35, 8'd3}: color_data = 12'h07a;
			{8'd35, 8'd4}: color_data = 12'h09d;
			{8'd35, 8'd5}: color_data = 12'h09d;
			{8'd35, 8'd6}: color_data = 12'h09d;
			{8'd35, 8'd7}: color_data = 12'h09d;
			{8'd35, 8'd8}: color_data = 12'h09d;
			{8'd35, 8'd9}: color_data = 12'h09d;
			{8'd35, 8'd10}: color_data = 12'h09d;
			{8'd35, 8'd11}: color_data = 12'h09d;
			{8'd35, 8'd12}: color_data = 12'h09d;
			{8'd35, 8'd13}: color_data = 12'h09d;
			{8'd35, 8'd14}: color_data = 12'h09d;
			{8'd35, 8'd15}: color_data = 12'h09d;
			{8'd35, 8'd16}: color_data = 12'h023;
			{8'd35, 8'd17}: color_data = 12'h000;
			{8'd35, 8'd18}: color_data = 12'h000;
			{8'd35, 8'd19}: color_data = 12'h000;
			{8'd35, 8'd20}: color_data = 12'h046;
			{8'd35, 8'd21}: color_data = 12'h0ad;
			{8'd35, 8'd22}: color_data = 12'h09d;
			{8'd35, 8'd23}: color_data = 12'h09d;
			{8'd35, 8'd24}: color_data = 12'h09d;
			{8'd35, 8'd25}: color_data = 12'h09d;
			{8'd35, 8'd26}: color_data = 12'h09d;
			{8'd35, 8'd27}: color_data = 12'h09d;
			{8'd35, 8'd28}: color_data = 12'h09d;
			{8'd35, 8'd29}: color_data = 12'h09d;
			{8'd35, 8'd30}: color_data = 12'h011;
			{8'd35, 8'd31}: color_data = 12'h000;
			{8'd35, 8'd32}: color_data = 12'h000;
			{8'd35, 8'd33}: color_data = 12'h000;
			{8'd35, 8'd34}: color_data = 12'h000;
			{8'd35, 8'd35}: color_data = 12'h000;
			{8'd35, 8'd36}: color_data = 12'h000;
			{8'd35, 8'd37}: color_data = 12'h000;
			{8'd35, 8'd38}: color_data = 12'h100;
			{8'd35, 8'd39}: color_data = 12'h710;
			{8'd35, 8'd40}: color_data = 12'hd20;
			{8'd35, 8'd41}: color_data = 12'hf21;
			{8'd35, 8'd42}: color_data = 12'he21;
			{8'd35, 8'd43}: color_data = 12'he21;
			{8'd35, 8'd44}: color_data = 12'he21;
			{8'd35, 8'd45}: color_data = 12'he21;
			{8'd35, 8'd46}: color_data = 12'he21;
			{8'd35, 8'd47}: color_data = 12'he21;
			{8'd35, 8'd48}: color_data = 12'he21;
			{8'd35, 8'd49}: color_data = 12'he21;
			{8'd35, 8'd50}: color_data = 12'he21;
			{8'd35, 8'd51}: color_data = 12'he21;
			{8'd35, 8'd52}: color_data = 12'he21;
			{8'd35, 8'd53}: color_data = 12'he21;
			{8'd35, 8'd54}: color_data = 12'h600;
			{8'd35, 8'd55}: color_data = 12'h000;
			{8'd35, 8'd56}: color_data = 12'h000;
			{8'd35, 8'd57}: color_data = 12'h000;
			{8'd35, 8'd58}: color_data = 12'h000;
			{8'd35, 8'd59}: color_data = 12'h000;
			{8'd35, 8'd60}: color_data = 12'h000;
			{8'd35, 8'd61}: color_data = 12'h000;
			{8'd35, 8'd62}: color_data = 12'h000;
			{8'd35, 8'd63}: color_data = 12'h000;
			{8'd35, 8'd100}: color_data = 12'he00;
			{8'd35, 8'd101}: color_data = 12'hf01;
			{8'd35, 8'd102}: color_data = 12'he00;
			{8'd35, 8'd103}: color_data = 12'he00;
			{8'd35, 8'd104}: color_data = 12'he00;
			{8'd35, 8'd105}: color_data = 12'he00;
			{8'd35, 8'd106}: color_data = 12'hc00;
			{8'd35, 8'd111}: color_data = 12'he01;
			{8'd35, 8'd112}: color_data = 12'he00;
			{8'd35, 8'd113}: color_data = 12'he00;
			{8'd35, 8'd114}: color_data = 12'he00;
			{8'd35, 8'd115}: color_data = 12'he00;
			{8'd35, 8'd116}: color_data = 12'he00;
			{8'd35, 8'd117}: color_data = 12'he00;
			{8'd35, 8'd118}: color_data = 12'he00;
			{8'd35, 8'd119}: color_data = 12'he00;
			{8'd35, 8'd120}: color_data = 12'he00;
			{8'd35, 8'd121}: color_data = 12'he00;
			{8'd35, 8'd122}: color_data = 12'he00;
			{8'd35, 8'd123}: color_data = 12'he00;
			{8'd35, 8'd124}: color_data = 12'he00;
			{8'd35, 8'd125}: color_data = 12'he00;
			{8'd35, 8'd126}: color_data = 12'he00;
			{8'd35, 8'd127}: color_data = 12'he00;
			{8'd35, 8'd128}: color_data = 12'he00;
			{8'd35, 8'd129}: color_data = 12'hb00;
			{8'd35, 8'd138}: color_data = 12'he00;
			{8'd35, 8'd139}: color_data = 12'he00;
			{8'd35, 8'd140}: color_data = 12'he00;
			{8'd35, 8'd141}: color_data = 12'he00;
			{8'd35, 8'd142}: color_data = 12'he00;
			{8'd35, 8'd143}: color_data = 12'he01;
			{8'd35, 8'd144}: color_data = 12'he00;
			{8'd36, 8'd0}: color_data = 12'h000;
			{8'd36, 8'd1}: color_data = 12'h000;
			{8'd36, 8'd2}: color_data = 12'h000;
			{8'd36, 8'd3}: color_data = 12'h08b;
			{8'd36, 8'd4}: color_data = 12'h09d;
			{8'd36, 8'd5}: color_data = 12'h09d;
			{8'd36, 8'd6}: color_data = 12'h09d;
			{8'd36, 8'd7}: color_data = 12'h09d;
			{8'd36, 8'd8}: color_data = 12'h09d;
			{8'd36, 8'd9}: color_data = 12'h09d;
			{8'd36, 8'd10}: color_data = 12'h09d;
			{8'd36, 8'd11}: color_data = 12'h09d;
			{8'd36, 8'd12}: color_data = 12'h09d;
			{8'd36, 8'd13}: color_data = 12'h09d;
			{8'd36, 8'd14}: color_data = 12'h09d;
			{8'd36, 8'd15}: color_data = 12'h0ae;
			{8'd36, 8'd16}: color_data = 12'h07a;
			{8'd36, 8'd17}: color_data = 12'h000;
			{8'd36, 8'd18}: color_data = 12'h000;
			{8'd36, 8'd19}: color_data = 12'h000;
			{8'd36, 8'd20}: color_data = 12'h000;
			{8'd36, 8'd21}: color_data = 12'h058;
			{8'd36, 8'd22}: color_data = 12'h0ae;
			{8'd36, 8'd23}: color_data = 12'h09d;
			{8'd36, 8'd24}: color_data = 12'h09d;
			{8'd36, 8'd25}: color_data = 12'h09d;
			{8'd36, 8'd26}: color_data = 12'h09d;
			{8'd36, 8'd27}: color_data = 12'h09d;
			{8'd36, 8'd28}: color_data = 12'h09d;
			{8'd36, 8'd29}: color_data = 12'h09d;
			{8'd36, 8'd30}: color_data = 12'h012;
			{8'd36, 8'd31}: color_data = 12'h000;
			{8'd36, 8'd32}: color_data = 12'h000;
			{8'd36, 8'd33}: color_data = 12'h000;
			{8'd36, 8'd34}: color_data = 12'h000;
			{8'd36, 8'd35}: color_data = 12'h000;
			{8'd36, 8'd36}: color_data = 12'h000;
			{8'd36, 8'd37}: color_data = 12'h610;
			{8'd36, 8'd38}: color_data = 12'hc10;
			{8'd36, 8'd39}: color_data = 12'he21;
			{8'd36, 8'd40}: color_data = 12'he21;
			{8'd36, 8'd41}: color_data = 12'he21;
			{8'd36, 8'd42}: color_data = 12'he21;
			{8'd36, 8'd43}: color_data = 12'he21;
			{8'd36, 8'd44}: color_data = 12'he21;
			{8'd36, 8'd45}: color_data = 12'he21;
			{8'd36, 8'd46}: color_data = 12'he21;
			{8'd36, 8'd47}: color_data = 12'he21;
			{8'd36, 8'd48}: color_data = 12'he21;
			{8'd36, 8'd49}: color_data = 12'he21;
			{8'd36, 8'd50}: color_data = 12'he21;
			{8'd36, 8'd51}: color_data = 12'he21;
			{8'd36, 8'd52}: color_data = 12'hd20;
			{8'd36, 8'd53}: color_data = 12'h400;
			{8'd36, 8'd54}: color_data = 12'h000;
			{8'd36, 8'd55}: color_data = 12'h000;
			{8'd36, 8'd56}: color_data = 12'h000;
			{8'd36, 8'd57}: color_data = 12'h000;
			{8'd36, 8'd58}: color_data = 12'h000;
			{8'd36, 8'd59}: color_data = 12'h000;
			{8'd36, 8'd60}: color_data = 12'h000;
			{8'd36, 8'd61}: color_data = 12'h000;
			{8'd36, 8'd62}: color_data = 12'h000;
			{8'd36, 8'd63}: color_data = 12'h000;
			{8'd36, 8'd64}: color_data = 12'h000;
			{8'd36, 8'd65}: color_data = 12'h000;
			{8'd36, 8'd66}: color_data = 12'h000;
			{8'd36, 8'd67}: color_data = 12'h000;
			{8'd36, 8'd68}: color_data = 12'h000;
			{8'd36, 8'd69}: color_data = 12'h000;
			{8'd36, 8'd70}: color_data = 12'h000;
			{8'd36, 8'd71}: color_data = 12'h000;
			{8'd36, 8'd72}: color_data = 12'h000;
			{8'd36, 8'd73}: color_data = 12'h000;
			{8'd36, 8'd74}: color_data = 12'h000;
			{8'd36, 8'd75}: color_data = 12'h000;
			{8'd36, 8'd100}: color_data = 12'he00;
			{8'd36, 8'd101}: color_data = 12'hf01;
			{8'd36, 8'd102}: color_data = 12'he00;
			{8'd36, 8'd103}: color_data = 12'he00;
			{8'd36, 8'd104}: color_data = 12'he00;
			{8'd36, 8'd105}: color_data = 12'he00;
			{8'd36, 8'd106}: color_data = 12'hc00;
			{8'd36, 8'd111}: color_data = 12'he00;
			{8'd36, 8'd112}: color_data = 12'he00;
			{8'd36, 8'd113}: color_data = 12'he00;
			{8'd36, 8'd114}: color_data = 12'he01;
			{8'd36, 8'd115}: color_data = 12'he01;
			{8'd36, 8'd116}: color_data = 12'he00;
			{8'd36, 8'd117}: color_data = 12'he00;
			{8'd36, 8'd118}: color_data = 12'he00;
			{8'd36, 8'd119}: color_data = 12'he00;
			{8'd36, 8'd120}: color_data = 12'he00;
			{8'd36, 8'd121}: color_data = 12'he00;
			{8'd36, 8'd122}: color_data = 12'he00;
			{8'd36, 8'd123}: color_data = 12'he00;
			{8'd36, 8'd124}: color_data = 12'he00;
			{8'd36, 8'd125}: color_data = 12'he00;
			{8'd36, 8'd126}: color_data = 12'he00;
			{8'd36, 8'd127}: color_data = 12'he01;
			{8'd36, 8'd128}: color_data = 12'he00;
			{8'd36, 8'd129}: color_data = 12'he00;
			{8'd36, 8'd130}: color_data = 12'he00;
			{8'd36, 8'd131}: color_data = 12'hd01;
			{8'd36, 8'd138}: color_data = 12'he00;
			{8'd36, 8'd139}: color_data = 12'he00;
			{8'd36, 8'd140}: color_data = 12'he00;
			{8'd36, 8'd141}: color_data = 12'he00;
			{8'd36, 8'd142}: color_data = 12'he00;
			{8'd36, 8'd143}: color_data = 12'he01;
			{8'd36, 8'd144}: color_data = 12'he00;
			{8'd37, 8'd0}: color_data = 12'h000;
			{8'd37, 8'd1}: color_data = 12'h000;
			{8'd37, 8'd2}: color_data = 12'h001;
			{8'd37, 8'd3}: color_data = 12'h08c;
			{8'd37, 8'd4}: color_data = 12'h09d;
			{8'd37, 8'd5}: color_data = 12'h09d;
			{8'd37, 8'd6}: color_data = 12'h09d;
			{8'd37, 8'd7}: color_data = 12'h09d;
			{8'd37, 8'd8}: color_data = 12'h09d;
			{8'd37, 8'd9}: color_data = 12'h09d;
			{8'd37, 8'd10}: color_data = 12'h09d;
			{8'd37, 8'd11}: color_data = 12'h09d;
			{8'd37, 8'd12}: color_data = 12'h09d;
			{8'd37, 8'd13}: color_data = 12'h09d;
			{8'd37, 8'd14}: color_data = 12'h09d;
			{8'd37, 8'd15}: color_data = 12'h09d;
			{8'd37, 8'd16}: color_data = 12'h0ae;
			{8'd37, 8'd17}: color_data = 12'h045;
			{8'd37, 8'd18}: color_data = 12'h000;
			{8'd37, 8'd19}: color_data = 12'h000;
			{8'd37, 8'd20}: color_data = 12'h000;
			{8'd37, 8'd21}: color_data = 12'h000;
			{8'd37, 8'd22}: color_data = 12'h069;
			{8'd37, 8'd23}: color_data = 12'h0ae;
			{8'd37, 8'd24}: color_data = 12'h09d;
			{8'd37, 8'd25}: color_data = 12'h09d;
			{8'd37, 8'd26}: color_data = 12'h09d;
			{8'd37, 8'd27}: color_data = 12'h09d;
			{8'd37, 8'd28}: color_data = 12'h09d;
			{8'd37, 8'd29}: color_data = 12'h09c;
			{8'd37, 8'd30}: color_data = 12'h011;
			{8'd37, 8'd31}: color_data = 12'h000;
			{8'd37, 8'd32}: color_data = 12'h000;
			{8'd37, 8'd33}: color_data = 12'h000;
			{8'd37, 8'd34}: color_data = 12'h000;
			{8'd37, 8'd35}: color_data = 12'h600;
			{8'd37, 8'd36}: color_data = 12'hc10;
			{8'd37, 8'd37}: color_data = 12'he21;
			{8'd37, 8'd38}: color_data = 12'he21;
			{8'd37, 8'd39}: color_data = 12'he21;
			{8'd37, 8'd40}: color_data = 12'he21;
			{8'd37, 8'd41}: color_data = 12'he21;
			{8'd37, 8'd42}: color_data = 12'he21;
			{8'd37, 8'd43}: color_data = 12'he21;
			{8'd37, 8'd44}: color_data = 12'he21;
			{8'd37, 8'd45}: color_data = 12'he21;
			{8'd37, 8'd46}: color_data = 12'he21;
			{8'd37, 8'd47}: color_data = 12'he21;
			{8'd37, 8'd48}: color_data = 12'he21;
			{8'd37, 8'd49}: color_data = 12'he21;
			{8'd37, 8'd50}: color_data = 12'he21;
			{8'd37, 8'd51}: color_data = 12'hb10;
			{8'd37, 8'd52}: color_data = 12'h100;
			{8'd37, 8'd53}: color_data = 12'h000;
			{8'd37, 8'd54}: color_data = 12'h000;
			{8'd37, 8'd55}: color_data = 12'h000;
			{8'd37, 8'd56}: color_data = 12'h000;
			{8'd37, 8'd57}: color_data = 12'h000;
			{8'd37, 8'd58}: color_data = 12'h000;
			{8'd37, 8'd59}: color_data = 12'h000;
			{8'd37, 8'd60}: color_data = 12'h000;
			{8'd37, 8'd61}: color_data = 12'h000;
			{8'd37, 8'd62}: color_data = 12'h000;
			{8'd37, 8'd63}: color_data = 12'h000;
			{8'd37, 8'd64}: color_data = 12'h000;
			{8'd37, 8'd65}: color_data = 12'h000;
			{8'd37, 8'd66}: color_data = 12'h000;
			{8'd37, 8'd67}: color_data = 12'h000;
			{8'd37, 8'd68}: color_data = 12'h000;
			{8'd37, 8'd69}: color_data = 12'h000;
			{8'd37, 8'd70}: color_data = 12'h000;
			{8'd37, 8'd71}: color_data = 12'h000;
			{8'd37, 8'd72}: color_data = 12'h000;
			{8'd37, 8'd73}: color_data = 12'h000;
			{8'd37, 8'd74}: color_data = 12'h000;
			{8'd37, 8'd75}: color_data = 12'h000;
			{8'd37, 8'd76}: color_data = 12'h000;
			{8'd37, 8'd100}: color_data = 12'he00;
			{8'd37, 8'd101}: color_data = 12'hf01;
			{8'd37, 8'd102}: color_data = 12'he00;
			{8'd37, 8'd103}: color_data = 12'he00;
			{8'd37, 8'd104}: color_data = 12'he00;
			{8'd37, 8'd105}: color_data = 12'he00;
			{8'd37, 8'd106}: color_data = 12'hc00;
			{8'd37, 8'd113}: color_data = 12'he01;
			{8'd37, 8'd114}: color_data = 12'he00;
			{8'd37, 8'd115}: color_data = 12'he00;
			{8'd37, 8'd116}: color_data = 12'he00;
			{8'd37, 8'd117}: color_data = 12'he00;
			{8'd37, 8'd118}: color_data = 12'he01;
			{8'd37, 8'd119}: color_data = 12'he00;
			{8'd37, 8'd120}: color_data = 12'he00;
			{8'd37, 8'd121}: color_data = 12'he00;
			{8'd37, 8'd122}: color_data = 12'he00;
			{8'd37, 8'd123}: color_data = 12'he00;
			{8'd37, 8'd124}: color_data = 12'he00;
			{8'd37, 8'd125}: color_data = 12'he00;
			{8'd37, 8'd126}: color_data = 12'he00;
			{8'd37, 8'd127}: color_data = 12'he00;
			{8'd37, 8'd128}: color_data = 12'he00;
			{8'd37, 8'd129}: color_data = 12'he00;
			{8'd37, 8'd130}: color_data = 12'he01;
			{8'd37, 8'd131}: color_data = 12'he00;
			{8'd37, 8'd132}: color_data = 12'he00;
			{8'd37, 8'd133}: color_data = 12'he00;
			{8'd37, 8'd138}: color_data = 12'he00;
			{8'd37, 8'd139}: color_data = 12'he00;
			{8'd37, 8'd140}: color_data = 12'he00;
			{8'd37, 8'd141}: color_data = 12'he00;
			{8'd37, 8'd142}: color_data = 12'he00;
			{8'd37, 8'd143}: color_data = 12'he01;
			{8'd37, 8'd144}: color_data = 12'he00;
			{8'd38, 8'd0}: color_data = 12'h000;
			{8'd38, 8'd1}: color_data = 12'h000;
			{8'd38, 8'd2}: color_data = 12'h012;
			{8'd38, 8'd3}: color_data = 12'h09d;
			{8'd38, 8'd4}: color_data = 12'h09d;
			{8'd38, 8'd5}: color_data = 12'h09d;
			{8'd38, 8'd6}: color_data = 12'h09d;
			{8'd38, 8'd7}: color_data = 12'h09d;
			{8'd38, 8'd8}: color_data = 12'h09d;
			{8'd38, 8'd9}: color_data = 12'h09d;
			{8'd38, 8'd10}: color_data = 12'h09d;
			{8'd38, 8'd11}: color_data = 12'h0ae;
			{8'd38, 8'd12}: color_data = 12'h09d;
			{8'd38, 8'd13}: color_data = 12'h09d;
			{8'd38, 8'd14}: color_data = 12'h09d;
			{8'd38, 8'd15}: color_data = 12'h09d;
			{8'd38, 8'd16}: color_data = 12'h09d;
			{8'd38, 8'd17}: color_data = 12'h08c;
			{8'd38, 8'd18}: color_data = 12'h011;
			{8'd38, 8'd19}: color_data = 12'h000;
			{8'd38, 8'd20}: color_data = 12'h000;
			{8'd38, 8'd21}: color_data = 12'h000;
			{8'd38, 8'd22}: color_data = 12'h001;
			{8'd38, 8'd23}: color_data = 12'h07a;
			{8'd38, 8'd24}: color_data = 12'h09d;
			{8'd38, 8'd25}: color_data = 12'h09d;
			{8'd38, 8'd26}: color_data = 12'h09d;
			{8'd38, 8'd27}: color_data = 12'h09d;
			{8'd38, 8'd28}: color_data = 12'h09d;
			{8'd38, 8'd29}: color_data = 12'h09c;
			{8'd38, 8'd30}: color_data = 12'h011;
			{8'd38, 8'd31}: color_data = 12'h000;
			{8'd38, 8'd32}: color_data = 12'h000;
			{8'd38, 8'd33}: color_data = 12'h000;
			{8'd38, 8'd34}: color_data = 12'h500;
			{8'd38, 8'd35}: color_data = 12'hf21;
			{8'd38, 8'd36}: color_data = 12'he21;
			{8'd38, 8'd37}: color_data = 12'he21;
			{8'd38, 8'd38}: color_data = 12'he21;
			{8'd38, 8'd39}: color_data = 12'he21;
			{8'd38, 8'd40}: color_data = 12'he21;
			{8'd38, 8'd41}: color_data = 12'he21;
			{8'd38, 8'd42}: color_data = 12'he21;
			{8'd38, 8'd43}: color_data = 12'he21;
			{8'd38, 8'd44}: color_data = 12'he21;
			{8'd38, 8'd45}: color_data = 12'he21;
			{8'd38, 8'd46}: color_data = 12'he21;
			{8'd38, 8'd47}: color_data = 12'he21;
			{8'd38, 8'd48}: color_data = 12'he21;
			{8'd38, 8'd49}: color_data = 12'he21;
			{8'd38, 8'd50}: color_data = 12'hd20;
			{8'd38, 8'd51}: color_data = 12'h710;
			{8'd38, 8'd52}: color_data = 12'h400;
			{8'd38, 8'd53}: color_data = 12'h400;
			{8'd38, 8'd54}: color_data = 12'h300;
			{8'd38, 8'd55}: color_data = 12'h200;
			{8'd38, 8'd56}: color_data = 12'h200;
			{8'd38, 8'd57}: color_data = 12'h100;
			{8'd38, 8'd58}: color_data = 12'h100;
			{8'd38, 8'd59}: color_data = 12'h000;
			{8'd38, 8'd60}: color_data = 12'h000;
			{8'd38, 8'd61}: color_data = 12'h000;
			{8'd38, 8'd62}: color_data = 12'h000;
			{8'd38, 8'd63}: color_data = 12'h000;
			{8'd38, 8'd64}: color_data = 12'h000;
			{8'd38, 8'd65}: color_data = 12'h000;
			{8'd38, 8'd66}: color_data = 12'h000;
			{8'd38, 8'd67}: color_data = 12'h000;
			{8'd38, 8'd68}: color_data = 12'h000;
			{8'd38, 8'd69}: color_data = 12'h000;
			{8'd38, 8'd70}: color_data = 12'h000;
			{8'd38, 8'd71}: color_data = 12'h000;
			{8'd38, 8'd72}: color_data = 12'h000;
			{8'd38, 8'd73}: color_data = 12'h000;
			{8'd38, 8'd74}: color_data = 12'h000;
			{8'd38, 8'd75}: color_data = 12'h000;
			{8'd38, 8'd76}: color_data = 12'h000;
			{8'd38, 8'd100}: color_data = 12'he00;
			{8'd38, 8'd101}: color_data = 12'hf01;
			{8'd38, 8'd102}: color_data = 12'he00;
			{8'd38, 8'd103}: color_data = 12'he00;
			{8'd38, 8'd104}: color_data = 12'he00;
			{8'd38, 8'd105}: color_data = 12'he00;
			{8'd38, 8'd106}: color_data = 12'hc00;
			{8'd38, 8'd116}: color_data = 12'he00;
			{8'd38, 8'd117}: color_data = 12'he00;
			{8'd38, 8'd118}: color_data = 12'he00;
			{8'd38, 8'd119}: color_data = 12'he00;
			{8'd38, 8'd120}: color_data = 12'he00;
			{8'd38, 8'd121}: color_data = 12'he01;
			{8'd38, 8'd122}: color_data = 12'he00;
			{8'd38, 8'd123}: color_data = 12'he00;
			{8'd38, 8'd124}: color_data = 12'he00;
			{8'd38, 8'd125}: color_data = 12'he00;
			{8'd38, 8'd126}: color_data = 12'he00;
			{8'd38, 8'd127}: color_data = 12'he00;
			{8'd38, 8'd128}: color_data = 12'he00;
			{8'd38, 8'd129}: color_data = 12'he00;
			{8'd38, 8'd130}: color_data = 12'he00;
			{8'd38, 8'd131}: color_data = 12'he00;
			{8'd38, 8'd132}: color_data = 12'hf01;
			{8'd38, 8'd133}: color_data = 12'he00;
			{8'd38, 8'd138}: color_data = 12'he00;
			{8'd38, 8'd139}: color_data = 12'he00;
			{8'd38, 8'd140}: color_data = 12'he00;
			{8'd38, 8'd141}: color_data = 12'he00;
			{8'd38, 8'd142}: color_data = 12'he00;
			{8'd38, 8'd143}: color_data = 12'he01;
			{8'd38, 8'd144}: color_data = 12'he00;
			{8'd39, 8'd0}: color_data = 12'h000;
			{8'd39, 8'd1}: color_data = 12'h000;
			{8'd39, 8'd2}: color_data = 12'h022;
			{8'd39, 8'd3}: color_data = 12'h09d;
			{8'd39, 8'd4}: color_data = 12'h09d;
			{8'd39, 8'd5}: color_data = 12'h09d;
			{8'd39, 8'd6}: color_data = 12'h09d;
			{8'd39, 8'd7}: color_data = 12'h09d;
			{8'd39, 8'd8}: color_data = 12'h09d;
			{8'd39, 8'd9}: color_data = 12'h0ae;
			{8'd39, 8'd10}: color_data = 12'h09d;
			{8'd39, 8'd11}: color_data = 12'h069;
			{8'd39, 8'd12}: color_data = 12'h09d;
			{8'd39, 8'd13}: color_data = 12'h09d;
			{8'd39, 8'd14}: color_data = 12'h09d;
			{8'd39, 8'd15}: color_data = 12'h09d;
			{8'd39, 8'd16}: color_data = 12'h09d;
			{8'd39, 8'd17}: color_data = 12'h0ae;
			{8'd39, 8'd18}: color_data = 12'h058;
			{8'd39, 8'd19}: color_data = 12'h000;
			{8'd39, 8'd20}: color_data = 12'h000;
			{8'd39, 8'd21}: color_data = 12'h000;
			{8'd39, 8'd22}: color_data = 12'h012;
			{8'd39, 8'd23}: color_data = 12'h07a;
			{8'd39, 8'd24}: color_data = 12'h09d;
			{8'd39, 8'd25}: color_data = 12'h09d;
			{8'd39, 8'd26}: color_data = 12'h09d;
			{8'd39, 8'd27}: color_data = 12'h09d;
			{8'd39, 8'd28}: color_data = 12'h09d;
			{8'd39, 8'd29}: color_data = 12'h09c;
			{8'd39, 8'd30}: color_data = 12'h011;
			{8'd39, 8'd31}: color_data = 12'h000;
			{8'd39, 8'd32}: color_data = 12'h000;
			{8'd39, 8'd33}: color_data = 12'h000;
			{8'd39, 8'd34}: color_data = 12'h400;
			{8'd39, 8'd35}: color_data = 12'he21;
			{8'd39, 8'd36}: color_data = 12'he21;
			{8'd39, 8'd37}: color_data = 12'he21;
			{8'd39, 8'd38}: color_data = 12'he21;
			{8'd39, 8'd39}: color_data = 12'he21;
			{8'd39, 8'd40}: color_data = 12'he21;
			{8'd39, 8'd41}: color_data = 12'he21;
			{8'd39, 8'd42}: color_data = 12'he21;
			{8'd39, 8'd43}: color_data = 12'he21;
			{8'd39, 8'd44}: color_data = 12'he21;
			{8'd39, 8'd45}: color_data = 12'he21;
			{8'd39, 8'd46}: color_data = 12'he21;
			{8'd39, 8'd47}: color_data = 12'he21;
			{8'd39, 8'd48}: color_data = 12'he21;
			{8'd39, 8'd49}: color_data = 12'he21;
			{8'd39, 8'd50}: color_data = 12'he21;
			{8'd39, 8'd51}: color_data = 12'he21;
			{8'd39, 8'd52}: color_data = 12'he21;
			{8'd39, 8'd53}: color_data = 12'he21;
			{8'd39, 8'd54}: color_data = 12'he21;
			{8'd39, 8'd55}: color_data = 12'he21;
			{8'd39, 8'd56}: color_data = 12'he20;
			{8'd39, 8'd57}: color_data = 12'hd20;
			{8'd39, 8'd58}: color_data = 12'hd20;
			{8'd39, 8'd59}: color_data = 12'hc10;
			{8'd39, 8'd60}: color_data = 12'hc10;
			{8'd39, 8'd61}: color_data = 12'hb10;
			{8'd39, 8'd62}: color_data = 12'ha10;
			{8'd39, 8'd63}: color_data = 12'ha10;
			{8'd39, 8'd64}: color_data = 12'h910;
			{8'd39, 8'd65}: color_data = 12'h810;
			{8'd39, 8'd66}: color_data = 12'h710;
			{8'd39, 8'd67}: color_data = 12'h610;
			{8'd39, 8'd68}: color_data = 12'h500;
			{8'd39, 8'd69}: color_data = 12'h000;
			{8'd39, 8'd70}: color_data = 12'h000;
			{8'd39, 8'd71}: color_data = 12'h000;
			{8'd39, 8'd72}: color_data = 12'h000;
			{8'd39, 8'd73}: color_data = 12'h000;
			{8'd39, 8'd74}: color_data = 12'h000;
			{8'd39, 8'd75}: color_data = 12'h000;
			{8'd39, 8'd76}: color_data = 12'h000;
			{8'd39, 8'd100}: color_data = 12'he00;
			{8'd39, 8'd101}: color_data = 12'hf01;
			{8'd39, 8'd102}: color_data = 12'he00;
			{8'd39, 8'd103}: color_data = 12'he00;
			{8'd39, 8'd104}: color_data = 12'he00;
			{8'd39, 8'd105}: color_data = 12'he00;
			{8'd39, 8'd106}: color_data = 12'hc00;
			{8'd39, 8'd119}: color_data = 12'he00;
			{8'd39, 8'd120}: color_data = 12'he00;
			{8'd39, 8'd121}: color_data = 12'he00;
			{8'd39, 8'd122}: color_data = 12'he00;
			{8'd39, 8'd123}: color_data = 12'he00;
			{8'd39, 8'd124}: color_data = 12'he01;
			{8'd39, 8'd125}: color_data = 12'he00;
			{8'd39, 8'd126}: color_data = 12'he00;
			{8'd39, 8'd127}: color_data = 12'he00;
			{8'd39, 8'd128}: color_data = 12'he00;
			{8'd39, 8'd129}: color_data = 12'he00;
			{8'd39, 8'd130}: color_data = 12'he00;
			{8'd39, 8'd131}: color_data = 12'he00;
			{8'd39, 8'd132}: color_data = 12'hf01;
			{8'd39, 8'd133}: color_data = 12'he00;
			{8'd39, 8'd138}: color_data = 12'he00;
			{8'd39, 8'd139}: color_data = 12'he00;
			{8'd39, 8'd140}: color_data = 12'he00;
			{8'd39, 8'd141}: color_data = 12'he00;
			{8'd39, 8'd142}: color_data = 12'he00;
			{8'd39, 8'd143}: color_data = 12'he01;
			{8'd39, 8'd144}: color_data = 12'he00;
			{8'd40, 8'd0}: color_data = 12'h000;
			{8'd40, 8'd1}: color_data = 12'h000;
			{8'd40, 8'd2}: color_data = 12'h024;
			{8'd40, 8'd3}: color_data = 12'h09d;
			{8'd40, 8'd4}: color_data = 12'h09d;
			{8'd40, 8'd5}: color_data = 12'h09d;
			{8'd40, 8'd6}: color_data = 12'h09d;
			{8'd40, 8'd7}: color_data = 12'h09d;
			{8'd40, 8'd8}: color_data = 12'h09d;
			{8'd40, 8'd9}: color_data = 12'h07a;
			{8'd40, 8'd10}: color_data = 12'h023;
			{8'd40, 8'd11}: color_data = 12'h000;
			{8'd40, 8'd12}: color_data = 12'h068;
			{8'd40, 8'd13}: color_data = 12'h0ae;
			{8'd40, 8'd14}: color_data = 12'h09d;
			{8'd40, 8'd15}: color_data = 12'h09d;
			{8'd40, 8'd16}: color_data = 12'h09d;
			{8'd40, 8'd17}: color_data = 12'h09d;
			{8'd40, 8'd18}: color_data = 12'h09d;
			{8'd40, 8'd19}: color_data = 12'h023;
			{8'd40, 8'd20}: color_data = 12'h000;
			{8'd40, 8'd21}: color_data = 12'h034;
			{8'd40, 8'd22}: color_data = 12'h09c;
			{8'd40, 8'd23}: color_data = 12'h09d;
			{8'd40, 8'd24}: color_data = 12'h09d;
			{8'd40, 8'd25}: color_data = 12'h09d;
			{8'd40, 8'd26}: color_data = 12'h09d;
			{8'd40, 8'd27}: color_data = 12'h09d;
			{8'd40, 8'd28}: color_data = 12'h09d;
			{8'd40, 8'd29}: color_data = 12'h09c;
			{8'd40, 8'd30}: color_data = 12'h001;
			{8'd40, 8'd31}: color_data = 12'h000;
			{8'd40, 8'd32}: color_data = 12'h000;
			{8'd40, 8'd33}: color_data = 12'h000;
			{8'd40, 8'd34}: color_data = 12'h200;
			{8'd40, 8'd35}: color_data = 12'he21;
			{8'd40, 8'd36}: color_data = 12'he21;
			{8'd40, 8'd37}: color_data = 12'he21;
			{8'd40, 8'd38}: color_data = 12'he21;
			{8'd40, 8'd39}: color_data = 12'he21;
			{8'd40, 8'd40}: color_data = 12'he21;
			{8'd40, 8'd41}: color_data = 12'he21;
			{8'd40, 8'd42}: color_data = 12'he21;
			{8'd40, 8'd43}: color_data = 12'he21;
			{8'd40, 8'd44}: color_data = 12'he21;
			{8'd40, 8'd45}: color_data = 12'he21;
			{8'd40, 8'd46}: color_data = 12'he21;
			{8'd40, 8'd47}: color_data = 12'he21;
			{8'd40, 8'd48}: color_data = 12'he21;
			{8'd40, 8'd49}: color_data = 12'he21;
			{8'd40, 8'd50}: color_data = 12'he21;
			{8'd40, 8'd51}: color_data = 12'he21;
			{8'd40, 8'd52}: color_data = 12'he21;
			{8'd40, 8'd53}: color_data = 12'he21;
			{8'd40, 8'd54}: color_data = 12'he21;
			{8'd40, 8'd55}: color_data = 12'he21;
			{8'd40, 8'd56}: color_data = 12'he21;
			{8'd40, 8'd57}: color_data = 12'he21;
			{8'd40, 8'd58}: color_data = 12'he21;
			{8'd40, 8'd59}: color_data = 12'he21;
			{8'd40, 8'd60}: color_data = 12'he21;
			{8'd40, 8'd61}: color_data = 12'he21;
			{8'd40, 8'd62}: color_data = 12'he21;
			{8'd40, 8'd63}: color_data = 12'he21;
			{8'd40, 8'd64}: color_data = 12'he21;
			{8'd40, 8'd65}: color_data = 12'he21;
			{8'd40, 8'd66}: color_data = 12'he21;
			{8'd40, 8'd67}: color_data = 12'hf21;
			{8'd40, 8'd68}: color_data = 12'he21;
			{8'd40, 8'd69}: color_data = 12'h200;
			{8'd40, 8'd70}: color_data = 12'h000;
			{8'd40, 8'd71}: color_data = 12'h000;
			{8'd40, 8'd72}: color_data = 12'h000;
			{8'd40, 8'd73}: color_data = 12'h000;
			{8'd40, 8'd74}: color_data = 12'h000;
			{8'd40, 8'd75}: color_data = 12'h000;
			{8'd40, 8'd76}: color_data = 12'h000;
			{8'd40, 8'd100}: color_data = 12'he00;
			{8'd40, 8'd101}: color_data = 12'hf01;
			{8'd40, 8'd102}: color_data = 12'he00;
			{8'd40, 8'd103}: color_data = 12'he00;
			{8'd40, 8'd104}: color_data = 12'he00;
			{8'd40, 8'd105}: color_data = 12'he00;
			{8'd40, 8'd106}: color_data = 12'hc00;
			{8'd40, 8'd122}: color_data = 12'he01;
			{8'd40, 8'd123}: color_data = 12'he01;
			{8'd40, 8'd124}: color_data = 12'he00;
			{8'd40, 8'd125}: color_data = 12'he00;
			{8'd40, 8'd126}: color_data = 12'he00;
			{8'd40, 8'd127}: color_data = 12'he00;
			{8'd40, 8'd128}: color_data = 12'he00;
			{8'd40, 8'd129}: color_data = 12'he00;
			{8'd40, 8'd130}: color_data = 12'he00;
			{8'd40, 8'd131}: color_data = 12'he00;
			{8'd40, 8'd132}: color_data = 12'hf01;
			{8'd40, 8'd133}: color_data = 12'he00;
			{8'd40, 8'd138}: color_data = 12'he00;
			{8'd40, 8'd139}: color_data = 12'he00;
			{8'd40, 8'd140}: color_data = 12'he00;
			{8'd40, 8'd141}: color_data = 12'he00;
			{8'd40, 8'd142}: color_data = 12'he00;
			{8'd40, 8'd143}: color_data = 12'he01;
			{8'd40, 8'd144}: color_data = 12'he00;
			{8'd41, 8'd0}: color_data = 12'h000;
			{8'd41, 8'd1}: color_data = 12'h000;
			{8'd41, 8'd2}: color_data = 12'h035;
			{8'd41, 8'd3}: color_data = 12'h0ae;
			{8'd41, 8'd4}: color_data = 12'h09d;
			{8'd41, 8'd5}: color_data = 12'h09d;
			{8'd41, 8'd6}: color_data = 12'h09d;
			{8'd41, 8'd7}: color_data = 12'h0ae;
			{8'd41, 8'd8}: color_data = 12'h068;
			{8'd41, 8'd9}: color_data = 12'h000;
			{8'd41, 8'd10}: color_data = 12'h000;
			{8'd41, 8'd11}: color_data = 12'h000;
			{8'd41, 8'd12}: color_data = 12'h001;
			{8'd41, 8'd13}: color_data = 12'h08b;
			{8'd41, 8'd14}: color_data = 12'h09d;
			{8'd41, 8'd15}: color_data = 12'h09d;
			{8'd41, 8'd16}: color_data = 12'h09d;
			{8'd41, 8'd17}: color_data = 12'h09d;
			{8'd41, 8'd18}: color_data = 12'h09d;
			{8'd41, 8'd19}: color_data = 12'h07a;
			{8'd41, 8'd20}: color_data = 12'h058;
			{8'd41, 8'd21}: color_data = 12'h09d;
			{8'd41, 8'd22}: color_data = 12'h09d;
			{8'd41, 8'd23}: color_data = 12'h09d;
			{8'd41, 8'd24}: color_data = 12'h09d;
			{8'd41, 8'd25}: color_data = 12'h09d;
			{8'd41, 8'd26}: color_data = 12'h09d;
			{8'd41, 8'd27}: color_data = 12'h09d;
			{8'd41, 8'd28}: color_data = 12'h09d;
			{8'd41, 8'd29}: color_data = 12'h08c;
			{8'd41, 8'd30}: color_data = 12'h001;
			{8'd41, 8'd31}: color_data = 12'h000;
			{8'd41, 8'd32}: color_data = 12'h000;
			{8'd41, 8'd33}: color_data = 12'h000;
			{8'd41, 8'd34}: color_data = 12'h100;
			{8'd41, 8'd35}: color_data = 12'hd20;
			{8'd41, 8'd36}: color_data = 12'he21;
			{8'd41, 8'd37}: color_data = 12'he21;
			{8'd41, 8'd38}: color_data = 12'he21;
			{8'd41, 8'd39}: color_data = 12'he21;
			{8'd41, 8'd40}: color_data = 12'he21;
			{8'd41, 8'd41}: color_data = 12'he21;
			{8'd41, 8'd42}: color_data = 12'he21;
			{8'd41, 8'd43}: color_data = 12'he21;
			{8'd41, 8'd44}: color_data = 12'he21;
			{8'd41, 8'd45}: color_data = 12'he21;
			{8'd41, 8'd46}: color_data = 12'he21;
			{8'd41, 8'd47}: color_data = 12'he21;
			{8'd41, 8'd48}: color_data = 12'he21;
			{8'd41, 8'd49}: color_data = 12'he21;
			{8'd41, 8'd50}: color_data = 12'he21;
			{8'd41, 8'd51}: color_data = 12'he21;
			{8'd41, 8'd52}: color_data = 12'he21;
			{8'd41, 8'd53}: color_data = 12'he21;
			{8'd41, 8'd54}: color_data = 12'he21;
			{8'd41, 8'd55}: color_data = 12'he21;
			{8'd41, 8'd56}: color_data = 12'he21;
			{8'd41, 8'd57}: color_data = 12'he21;
			{8'd41, 8'd58}: color_data = 12'he21;
			{8'd41, 8'd59}: color_data = 12'he21;
			{8'd41, 8'd60}: color_data = 12'he21;
			{8'd41, 8'd61}: color_data = 12'he21;
			{8'd41, 8'd62}: color_data = 12'he21;
			{8'd41, 8'd63}: color_data = 12'he21;
			{8'd41, 8'd64}: color_data = 12'he21;
			{8'd41, 8'd65}: color_data = 12'he21;
			{8'd41, 8'd66}: color_data = 12'he21;
			{8'd41, 8'd67}: color_data = 12'he21;
			{8'd41, 8'd68}: color_data = 12'hc10;
			{8'd41, 8'd69}: color_data = 12'h000;
			{8'd41, 8'd70}: color_data = 12'h000;
			{8'd41, 8'd71}: color_data = 12'h000;
			{8'd41, 8'd72}: color_data = 12'h000;
			{8'd41, 8'd73}: color_data = 12'h000;
			{8'd41, 8'd74}: color_data = 12'h000;
			{8'd41, 8'd75}: color_data = 12'h000;
			{8'd41, 8'd100}: color_data = 12'he00;
			{8'd41, 8'd101}: color_data = 12'hf01;
			{8'd41, 8'd102}: color_data = 12'he00;
			{8'd41, 8'd103}: color_data = 12'he00;
			{8'd41, 8'd104}: color_data = 12'he00;
			{8'd41, 8'd105}: color_data = 12'he00;
			{8'd41, 8'd106}: color_data = 12'hc00;
			{8'd41, 8'd125}: color_data = 12'he00;
			{8'd41, 8'd126}: color_data = 12'he00;
			{8'd41, 8'd127}: color_data = 12'he00;
			{8'd41, 8'd128}: color_data = 12'he00;
			{8'd41, 8'd129}: color_data = 12'he00;
			{8'd41, 8'd130}: color_data = 12'he00;
			{8'd41, 8'd131}: color_data = 12'he00;
			{8'd41, 8'd132}: color_data = 12'hf01;
			{8'd41, 8'd133}: color_data = 12'he00;
			{8'd41, 8'd138}: color_data = 12'he00;
			{8'd41, 8'd139}: color_data = 12'he00;
			{8'd41, 8'd140}: color_data = 12'he00;
			{8'd41, 8'd141}: color_data = 12'he00;
			{8'd41, 8'd142}: color_data = 12'he00;
			{8'd41, 8'd143}: color_data = 12'he01;
			{8'd41, 8'd144}: color_data = 12'he00;
			{8'd42, 8'd0}: color_data = 12'h000;
			{8'd42, 8'd1}: color_data = 12'h000;
			{8'd42, 8'd2}: color_data = 12'h046;
			{8'd42, 8'd3}: color_data = 12'h0ae;
			{8'd42, 8'd4}: color_data = 12'h09d;
			{8'd42, 8'd5}: color_data = 12'h09d;
			{8'd42, 8'd6}: color_data = 12'h09d;
			{8'd42, 8'd7}: color_data = 12'h09d;
			{8'd42, 8'd8}: color_data = 12'h08b;
			{8'd42, 8'd9}: color_data = 12'h011;
			{8'd42, 8'd10}: color_data = 12'h000;
			{8'd42, 8'd11}: color_data = 12'h000;
			{8'd42, 8'd12}: color_data = 12'h000;
			{8'd42, 8'd13}: color_data = 12'h034;
			{8'd42, 8'd14}: color_data = 12'h09d;
			{8'd42, 8'd15}: color_data = 12'h09d;
			{8'd42, 8'd16}: color_data = 12'h09d;
			{8'd42, 8'd17}: color_data = 12'h09d;
			{8'd42, 8'd18}: color_data = 12'h09d;
			{8'd42, 8'd19}: color_data = 12'h09d;
			{8'd42, 8'd20}: color_data = 12'h0ae;
			{8'd42, 8'd21}: color_data = 12'h09d;
			{8'd42, 8'd22}: color_data = 12'h09d;
			{8'd42, 8'd23}: color_data = 12'h09d;
			{8'd42, 8'd24}: color_data = 12'h09d;
			{8'd42, 8'd25}: color_data = 12'h09d;
			{8'd42, 8'd26}: color_data = 12'h09d;
			{8'd42, 8'd27}: color_data = 12'h09d;
			{8'd42, 8'd28}: color_data = 12'h09d;
			{8'd42, 8'd29}: color_data = 12'h08c;
			{8'd42, 8'd30}: color_data = 12'h001;
			{8'd42, 8'd31}: color_data = 12'h000;
			{8'd42, 8'd32}: color_data = 12'h000;
			{8'd42, 8'd33}: color_data = 12'h000;
			{8'd42, 8'd34}: color_data = 12'h000;
			{8'd42, 8'd35}: color_data = 12'hc10;
			{8'd42, 8'd36}: color_data = 12'he21;
			{8'd42, 8'd37}: color_data = 12'he21;
			{8'd42, 8'd38}: color_data = 12'he21;
			{8'd42, 8'd39}: color_data = 12'he21;
			{8'd42, 8'd40}: color_data = 12'he21;
			{8'd42, 8'd41}: color_data = 12'he21;
			{8'd42, 8'd42}: color_data = 12'he21;
			{8'd42, 8'd43}: color_data = 12'he21;
			{8'd42, 8'd44}: color_data = 12'he21;
			{8'd42, 8'd45}: color_data = 12'he21;
			{8'd42, 8'd46}: color_data = 12'he21;
			{8'd42, 8'd47}: color_data = 12'he21;
			{8'd42, 8'd48}: color_data = 12'he21;
			{8'd42, 8'd49}: color_data = 12'he21;
			{8'd42, 8'd50}: color_data = 12'he21;
			{8'd42, 8'd51}: color_data = 12'he21;
			{8'd42, 8'd52}: color_data = 12'he21;
			{8'd42, 8'd53}: color_data = 12'he21;
			{8'd42, 8'd54}: color_data = 12'he21;
			{8'd42, 8'd55}: color_data = 12'he21;
			{8'd42, 8'd56}: color_data = 12'he21;
			{8'd42, 8'd57}: color_data = 12'he21;
			{8'd42, 8'd58}: color_data = 12'he21;
			{8'd42, 8'd59}: color_data = 12'he21;
			{8'd42, 8'd60}: color_data = 12'he21;
			{8'd42, 8'd61}: color_data = 12'he21;
			{8'd42, 8'd62}: color_data = 12'he21;
			{8'd42, 8'd63}: color_data = 12'he21;
			{8'd42, 8'd64}: color_data = 12'he21;
			{8'd42, 8'd65}: color_data = 12'he21;
			{8'd42, 8'd66}: color_data = 12'he21;
			{8'd42, 8'd67}: color_data = 12'he21;
			{8'd42, 8'd68}: color_data = 12'h910;
			{8'd42, 8'd69}: color_data = 12'h000;
			{8'd42, 8'd70}: color_data = 12'h000;
			{8'd42, 8'd71}: color_data = 12'h000;
			{8'd42, 8'd72}: color_data = 12'h000;
			{8'd42, 8'd73}: color_data = 12'h000;
			{8'd42, 8'd74}: color_data = 12'h000;
			{8'd42, 8'd75}: color_data = 12'h000;
			{8'd42, 8'd100}: color_data = 12'he00;
			{8'd42, 8'd101}: color_data = 12'hf01;
			{8'd42, 8'd102}: color_data = 12'he00;
			{8'd42, 8'd103}: color_data = 12'he00;
			{8'd42, 8'd104}: color_data = 12'he00;
			{8'd42, 8'd105}: color_data = 12'he00;
			{8'd42, 8'd106}: color_data = 12'hc00;
			{8'd42, 8'd121}: color_data = 12'hf00;
			{8'd42, 8'd122}: color_data = 12'he00;
			{8'd42, 8'd123}: color_data = 12'he00;
			{8'd42, 8'd124}: color_data = 12'he01;
			{8'd42, 8'd125}: color_data = 12'he00;
			{8'd42, 8'd126}: color_data = 12'he00;
			{8'd42, 8'd127}: color_data = 12'he00;
			{8'd42, 8'd128}: color_data = 12'he00;
			{8'd42, 8'd129}: color_data = 12'he00;
			{8'd42, 8'd130}: color_data = 12'he00;
			{8'd42, 8'd131}: color_data = 12'he00;
			{8'd42, 8'd132}: color_data = 12'hf01;
			{8'd42, 8'd133}: color_data = 12'he00;
			{8'd42, 8'd138}: color_data = 12'he00;
			{8'd42, 8'd139}: color_data = 12'he00;
			{8'd42, 8'd140}: color_data = 12'he00;
			{8'd42, 8'd141}: color_data = 12'he00;
			{8'd42, 8'd142}: color_data = 12'he00;
			{8'd42, 8'd143}: color_data = 12'he01;
			{8'd42, 8'd144}: color_data = 12'he00;
			{8'd43, 8'd0}: color_data = 12'h000;
			{8'd43, 8'd1}: color_data = 12'h000;
			{8'd43, 8'd2}: color_data = 12'h057;
			{8'd43, 8'd3}: color_data = 12'h0ae;
			{8'd43, 8'd4}: color_data = 12'h09d;
			{8'd43, 8'd5}: color_data = 12'h09d;
			{8'd43, 8'd6}: color_data = 12'h09d;
			{8'd43, 8'd7}: color_data = 12'h09d;
			{8'd43, 8'd8}: color_data = 12'h0ae;
			{8'd43, 8'd9}: color_data = 12'h068;
			{8'd43, 8'd10}: color_data = 12'h000;
			{8'd43, 8'd11}: color_data = 12'h000;
			{8'd43, 8'd12}: color_data = 12'h000;
			{8'd43, 8'd13}: color_data = 12'h000;
			{8'd43, 8'd14}: color_data = 12'h068;
			{8'd43, 8'd15}: color_data = 12'h0ae;
			{8'd43, 8'd16}: color_data = 12'h09d;
			{8'd43, 8'd17}: color_data = 12'h09d;
			{8'd43, 8'd18}: color_data = 12'h09d;
			{8'd43, 8'd19}: color_data = 12'h09d;
			{8'd43, 8'd20}: color_data = 12'h09d;
			{8'd43, 8'd21}: color_data = 12'h09d;
			{8'd43, 8'd22}: color_data = 12'h09d;
			{8'd43, 8'd23}: color_data = 12'h09d;
			{8'd43, 8'd24}: color_data = 12'h09d;
			{8'd43, 8'd25}: color_data = 12'h09d;
			{8'd43, 8'd26}: color_data = 12'h09d;
			{8'd43, 8'd27}: color_data = 12'h09d;
			{8'd43, 8'd28}: color_data = 12'h09d;
			{8'd43, 8'd29}: color_data = 12'h08c;
			{8'd43, 8'd30}: color_data = 12'h000;
			{8'd43, 8'd31}: color_data = 12'h000;
			{8'd43, 8'd32}: color_data = 12'h000;
			{8'd43, 8'd33}: color_data = 12'h000;
			{8'd43, 8'd34}: color_data = 12'h000;
			{8'd43, 8'd35}: color_data = 12'ha10;
			{8'd43, 8'd36}: color_data = 12'he21;
			{8'd43, 8'd37}: color_data = 12'he21;
			{8'd43, 8'd38}: color_data = 12'he21;
			{8'd43, 8'd39}: color_data = 12'he21;
			{8'd43, 8'd40}: color_data = 12'he21;
			{8'd43, 8'd41}: color_data = 12'he21;
			{8'd43, 8'd42}: color_data = 12'he21;
			{8'd43, 8'd43}: color_data = 12'he21;
			{8'd43, 8'd44}: color_data = 12'he21;
			{8'd43, 8'd45}: color_data = 12'he21;
			{8'd43, 8'd46}: color_data = 12'he21;
			{8'd43, 8'd47}: color_data = 12'he21;
			{8'd43, 8'd48}: color_data = 12'he21;
			{8'd43, 8'd49}: color_data = 12'he21;
			{8'd43, 8'd50}: color_data = 12'he21;
			{8'd43, 8'd51}: color_data = 12'he21;
			{8'd43, 8'd52}: color_data = 12'he21;
			{8'd43, 8'd53}: color_data = 12'he21;
			{8'd43, 8'd54}: color_data = 12'he21;
			{8'd43, 8'd55}: color_data = 12'he21;
			{8'd43, 8'd56}: color_data = 12'he21;
			{8'd43, 8'd57}: color_data = 12'he21;
			{8'd43, 8'd58}: color_data = 12'he21;
			{8'd43, 8'd59}: color_data = 12'he21;
			{8'd43, 8'd60}: color_data = 12'he21;
			{8'd43, 8'd61}: color_data = 12'he21;
			{8'd43, 8'd62}: color_data = 12'he21;
			{8'd43, 8'd63}: color_data = 12'he21;
			{8'd43, 8'd64}: color_data = 12'he21;
			{8'd43, 8'd65}: color_data = 12'he21;
			{8'd43, 8'd66}: color_data = 12'he21;
			{8'd43, 8'd67}: color_data = 12'he21;
			{8'd43, 8'd68}: color_data = 12'h610;
			{8'd43, 8'd69}: color_data = 12'h000;
			{8'd43, 8'd70}: color_data = 12'h000;
			{8'd43, 8'd71}: color_data = 12'h000;
			{8'd43, 8'd72}: color_data = 12'h000;
			{8'd43, 8'd73}: color_data = 12'h000;
			{8'd43, 8'd74}: color_data = 12'h000;
			{8'd43, 8'd75}: color_data = 12'h000;
			{8'd43, 8'd100}: color_data = 12'he00;
			{8'd43, 8'd101}: color_data = 12'hf01;
			{8'd43, 8'd102}: color_data = 12'he00;
			{8'd43, 8'd103}: color_data = 12'he00;
			{8'd43, 8'd104}: color_data = 12'he00;
			{8'd43, 8'd105}: color_data = 12'he00;
			{8'd43, 8'd106}: color_data = 12'hc00;
			{8'd43, 8'd118}: color_data = 12'hf00;
			{8'd43, 8'd119}: color_data = 12'he00;
			{8'd43, 8'd120}: color_data = 12'he00;
			{8'd43, 8'd121}: color_data = 12'he00;
			{8'd43, 8'd122}: color_data = 12'he00;
			{8'd43, 8'd123}: color_data = 12'he01;
			{8'd43, 8'd124}: color_data = 12'he01;
			{8'd43, 8'd125}: color_data = 12'he00;
			{8'd43, 8'd126}: color_data = 12'he00;
			{8'd43, 8'd127}: color_data = 12'he00;
			{8'd43, 8'd128}: color_data = 12'he00;
			{8'd43, 8'd129}: color_data = 12'he00;
			{8'd43, 8'd130}: color_data = 12'he00;
			{8'd43, 8'd131}: color_data = 12'he00;
			{8'd43, 8'd132}: color_data = 12'hf01;
			{8'd43, 8'd133}: color_data = 12'he00;
			{8'd43, 8'd138}: color_data = 12'he00;
			{8'd43, 8'd139}: color_data = 12'he00;
			{8'd43, 8'd140}: color_data = 12'he00;
			{8'd43, 8'd141}: color_data = 12'he00;
			{8'd43, 8'd142}: color_data = 12'he00;
			{8'd43, 8'd143}: color_data = 12'he01;
			{8'd43, 8'd144}: color_data = 12'he00;
			{8'd44, 8'd0}: color_data = 12'h000;
			{8'd44, 8'd1}: color_data = 12'h000;
			{8'd44, 8'd2}: color_data = 12'h069;
			{8'd44, 8'd3}: color_data = 12'h0ae;
			{8'd44, 8'd4}: color_data = 12'h09d;
			{8'd44, 8'd5}: color_data = 12'h09d;
			{8'd44, 8'd6}: color_data = 12'h09d;
			{8'd44, 8'd7}: color_data = 12'h09d;
			{8'd44, 8'd8}: color_data = 12'h09d;
			{8'd44, 8'd9}: color_data = 12'h09d;
			{8'd44, 8'd10}: color_data = 12'h035;
			{8'd44, 8'd11}: color_data = 12'h000;
			{8'd44, 8'd12}: color_data = 12'h000;
			{8'd44, 8'd13}: color_data = 12'h000;
			{8'd44, 8'd14}: color_data = 12'h011;
			{8'd44, 8'd15}: color_data = 12'h08c;
			{8'd44, 8'd16}: color_data = 12'h09d;
			{8'd44, 8'd17}: color_data = 12'h09d;
			{8'd44, 8'd18}: color_data = 12'h09d;
			{8'd44, 8'd19}: color_data = 12'h09d;
			{8'd44, 8'd20}: color_data = 12'h09d;
			{8'd44, 8'd21}: color_data = 12'h09d;
			{8'd44, 8'd22}: color_data = 12'h09d;
			{8'd44, 8'd23}: color_data = 12'h09d;
			{8'd44, 8'd24}: color_data = 12'h09d;
			{8'd44, 8'd25}: color_data = 12'h09d;
			{8'd44, 8'd26}: color_data = 12'h09d;
			{8'd44, 8'd27}: color_data = 12'h09d;
			{8'd44, 8'd28}: color_data = 12'h09d;
			{8'd44, 8'd29}: color_data = 12'h08c;
			{8'd44, 8'd30}: color_data = 12'h000;
			{8'd44, 8'd31}: color_data = 12'h000;
			{8'd44, 8'd32}: color_data = 12'h000;
			{8'd44, 8'd33}: color_data = 12'h000;
			{8'd44, 8'd34}: color_data = 12'h000;
			{8'd44, 8'd35}: color_data = 12'h810;
			{8'd44, 8'd36}: color_data = 12'he21;
			{8'd44, 8'd37}: color_data = 12'he21;
			{8'd44, 8'd38}: color_data = 12'he21;
			{8'd44, 8'd39}: color_data = 12'he21;
			{8'd44, 8'd40}: color_data = 12'he21;
			{8'd44, 8'd41}: color_data = 12'he21;
			{8'd44, 8'd42}: color_data = 12'he21;
			{8'd44, 8'd43}: color_data = 12'he21;
			{8'd44, 8'd44}: color_data = 12'he21;
			{8'd44, 8'd45}: color_data = 12'he21;
			{8'd44, 8'd46}: color_data = 12'he21;
			{8'd44, 8'd47}: color_data = 12'he21;
			{8'd44, 8'd48}: color_data = 12'he21;
			{8'd44, 8'd49}: color_data = 12'he21;
			{8'd44, 8'd50}: color_data = 12'he21;
			{8'd44, 8'd51}: color_data = 12'he21;
			{8'd44, 8'd52}: color_data = 12'he21;
			{8'd44, 8'd53}: color_data = 12'he21;
			{8'd44, 8'd54}: color_data = 12'he21;
			{8'd44, 8'd55}: color_data = 12'he21;
			{8'd44, 8'd56}: color_data = 12'he21;
			{8'd44, 8'd57}: color_data = 12'he21;
			{8'd44, 8'd58}: color_data = 12'he21;
			{8'd44, 8'd59}: color_data = 12'he21;
			{8'd44, 8'd60}: color_data = 12'he21;
			{8'd44, 8'd61}: color_data = 12'he21;
			{8'd44, 8'd62}: color_data = 12'he21;
			{8'd44, 8'd63}: color_data = 12'he21;
			{8'd44, 8'd64}: color_data = 12'he21;
			{8'd44, 8'd65}: color_data = 12'he21;
			{8'd44, 8'd66}: color_data = 12'he21;
			{8'd44, 8'd67}: color_data = 12'he21;
			{8'd44, 8'd68}: color_data = 12'h400;
			{8'd44, 8'd69}: color_data = 12'h000;
			{8'd44, 8'd70}: color_data = 12'h000;
			{8'd44, 8'd71}: color_data = 12'h000;
			{8'd44, 8'd72}: color_data = 12'h000;
			{8'd44, 8'd73}: color_data = 12'h000;
			{8'd44, 8'd74}: color_data = 12'h000;
			{8'd44, 8'd75}: color_data = 12'h000;
			{8'd44, 8'd100}: color_data = 12'he00;
			{8'd44, 8'd101}: color_data = 12'hf01;
			{8'd44, 8'd102}: color_data = 12'he00;
			{8'd44, 8'd103}: color_data = 12'he00;
			{8'd44, 8'd104}: color_data = 12'he00;
			{8'd44, 8'd105}: color_data = 12'he00;
			{8'd44, 8'd106}: color_data = 12'hc00;
			{8'd44, 8'd115}: color_data = 12'he01;
			{8'd44, 8'd116}: color_data = 12'he00;
			{8'd44, 8'd117}: color_data = 12'he00;
			{8'd44, 8'd118}: color_data = 12'he00;
			{8'd44, 8'd119}: color_data = 12'he00;
			{8'd44, 8'd120}: color_data = 12'he01;
			{8'd44, 8'd121}: color_data = 12'he00;
			{8'd44, 8'd122}: color_data = 12'he00;
			{8'd44, 8'd123}: color_data = 12'he00;
			{8'd44, 8'd124}: color_data = 12'he00;
			{8'd44, 8'd125}: color_data = 12'he00;
			{8'd44, 8'd126}: color_data = 12'he00;
			{8'd44, 8'd127}: color_data = 12'he00;
			{8'd44, 8'd128}: color_data = 12'he00;
			{8'd44, 8'd129}: color_data = 12'he00;
			{8'd44, 8'd130}: color_data = 12'he00;
			{8'd44, 8'd131}: color_data = 12'he00;
			{8'd44, 8'd132}: color_data = 12'hf01;
			{8'd44, 8'd133}: color_data = 12'he00;
			{8'd44, 8'd138}: color_data = 12'he00;
			{8'd44, 8'd139}: color_data = 12'he00;
			{8'd44, 8'd140}: color_data = 12'he00;
			{8'd44, 8'd141}: color_data = 12'he00;
			{8'd44, 8'd142}: color_data = 12'he00;
			{8'd44, 8'd143}: color_data = 12'he01;
			{8'd44, 8'd144}: color_data = 12'he00;
			{8'd45, 8'd0}: color_data = 12'h000;
			{8'd45, 8'd1}: color_data = 12'h000;
			{8'd45, 8'd2}: color_data = 12'h034;
			{8'd45, 8'd3}: color_data = 12'h09d;
			{8'd45, 8'd4}: color_data = 12'h09d;
			{8'd45, 8'd5}: color_data = 12'h09d;
			{8'd45, 8'd6}: color_data = 12'h09d;
			{8'd45, 8'd7}: color_data = 12'h09d;
			{8'd45, 8'd8}: color_data = 12'h09d;
			{8'd45, 8'd9}: color_data = 12'h09d;
			{8'd45, 8'd10}: color_data = 12'h08c;
			{8'd45, 8'd11}: color_data = 12'h011;
			{8'd45, 8'd12}: color_data = 12'h000;
			{8'd45, 8'd13}: color_data = 12'h000;
			{8'd45, 8'd14}: color_data = 12'h000;
			{8'd45, 8'd15}: color_data = 12'h034;
			{8'd45, 8'd16}: color_data = 12'h09d;
			{8'd45, 8'd17}: color_data = 12'h09d;
			{8'd45, 8'd18}: color_data = 12'h09d;
			{8'd45, 8'd19}: color_data = 12'h09d;
			{8'd45, 8'd20}: color_data = 12'h09d;
			{8'd45, 8'd21}: color_data = 12'h09d;
			{8'd45, 8'd22}: color_data = 12'h09d;
			{8'd45, 8'd23}: color_data = 12'h09d;
			{8'd45, 8'd24}: color_data = 12'h09d;
			{8'd45, 8'd25}: color_data = 12'h09d;
			{8'd45, 8'd26}: color_data = 12'h09d;
			{8'd45, 8'd27}: color_data = 12'h09d;
			{8'd45, 8'd28}: color_data = 12'h09d;
			{8'd45, 8'd29}: color_data = 12'h08b;
			{8'd45, 8'd30}: color_data = 12'h000;
			{8'd45, 8'd31}: color_data = 12'h000;
			{8'd45, 8'd32}: color_data = 12'h000;
			{8'd45, 8'd33}: color_data = 12'h000;
			{8'd45, 8'd34}: color_data = 12'h000;
			{8'd45, 8'd35}: color_data = 12'h710;
			{8'd45, 8'd36}: color_data = 12'hf21;
			{8'd45, 8'd37}: color_data = 12'he21;
			{8'd45, 8'd38}: color_data = 12'he21;
			{8'd45, 8'd39}: color_data = 12'he21;
			{8'd45, 8'd40}: color_data = 12'he21;
			{8'd45, 8'd41}: color_data = 12'he21;
			{8'd45, 8'd42}: color_data = 12'he21;
			{8'd45, 8'd43}: color_data = 12'he21;
			{8'd45, 8'd44}: color_data = 12'he21;
			{8'd45, 8'd45}: color_data = 12'he21;
			{8'd45, 8'd46}: color_data = 12'he21;
			{8'd45, 8'd47}: color_data = 12'he21;
			{8'd45, 8'd48}: color_data = 12'he21;
			{8'd45, 8'd49}: color_data = 12'he21;
			{8'd45, 8'd50}: color_data = 12'he21;
			{8'd45, 8'd51}: color_data = 12'he21;
			{8'd45, 8'd52}: color_data = 12'he21;
			{8'd45, 8'd53}: color_data = 12'he21;
			{8'd45, 8'd54}: color_data = 12'he21;
			{8'd45, 8'd55}: color_data = 12'he21;
			{8'd45, 8'd56}: color_data = 12'he21;
			{8'd45, 8'd57}: color_data = 12'he21;
			{8'd45, 8'd58}: color_data = 12'he21;
			{8'd45, 8'd59}: color_data = 12'he21;
			{8'd45, 8'd60}: color_data = 12'he21;
			{8'd45, 8'd61}: color_data = 12'he21;
			{8'd45, 8'd62}: color_data = 12'he21;
			{8'd45, 8'd63}: color_data = 12'he21;
			{8'd45, 8'd64}: color_data = 12'he21;
			{8'd45, 8'd65}: color_data = 12'he21;
			{8'd45, 8'd66}: color_data = 12'he21;
			{8'd45, 8'd67}: color_data = 12'hd20;
			{8'd45, 8'd68}: color_data = 12'h100;
			{8'd45, 8'd69}: color_data = 12'h000;
			{8'd45, 8'd70}: color_data = 12'h000;
			{8'd45, 8'd71}: color_data = 12'h000;
			{8'd45, 8'd72}: color_data = 12'h000;
			{8'd45, 8'd73}: color_data = 12'h000;
			{8'd45, 8'd74}: color_data = 12'h000;
			{8'd45, 8'd75}: color_data = 12'h000;
			{8'd45, 8'd100}: color_data = 12'he00;
			{8'd45, 8'd101}: color_data = 12'hf01;
			{8'd45, 8'd102}: color_data = 12'he00;
			{8'd45, 8'd103}: color_data = 12'he00;
			{8'd45, 8'd104}: color_data = 12'he00;
			{8'd45, 8'd105}: color_data = 12'he00;
			{8'd45, 8'd106}: color_data = 12'hc00;
			{8'd45, 8'd112}: color_data = 12'he00;
			{8'd45, 8'd113}: color_data = 12'he00;
			{8'd45, 8'd114}: color_data = 12'he00;
			{8'd45, 8'd115}: color_data = 12'he00;
			{8'd45, 8'd116}: color_data = 12'he00;
			{8'd45, 8'd117}: color_data = 12'he01;
			{8'd45, 8'd118}: color_data = 12'he00;
			{8'd45, 8'd119}: color_data = 12'he00;
			{8'd45, 8'd120}: color_data = 12'he00;
			{8'd45, 8'd121}: color_data = 12'he00;
			{8'd45, 8'd122}: color_data = 12'he00;
			{8'd45, 8'd123}: color_data = 12'he00;
			{8'd45, 8'd124}: color_data = 12'he00;
			{8'd45, 8'd125}: color_data = 12'he00;
			{8'd45, 8'd126}: color_data = 12'he00;
			{8'd45, 8'd127}: color_data = 12'he00;
			{8'd45, 8'd128}: color_data = 12'he00;
			{8'd45, 8'd129}: color_data = 12'hf01;
			{8'd45, 8'd130}: color_data = 12'he00;
			{8'd45, 8'd131}: color_data = 12'he00;
			{8'd45, 8'd132}: color_data = 12'he00;
			{8'd45, 8'd133}: color_data = 12'he00;
			{8'd45, 8'd138}: color_data = 12'he00;
			{8'd45, 8'd139}: color_data = 12'he00;
			{8'd45, 8'd140}: color_data = 12'he00;
			{8'd45, 8'd141}: color_data = 12'he00;
			{8'd45, 8'd142}: color_data = 12'he00;
			{8'd45, 8'd143}: color_data = 12'he01;
			{8'd45, 8'd144}: color_data = 12'he00;
			{8'd46, 8'd0}: color_data = 12'h000;
			{8'd46, 8'd1}: color_data = 12'h000;
			{8'd46, 8'd2}: color_data = 12'h000;
			{8'd46, 8'd3}: color_data = 12'h057;
			{8'd46, 8'd4}: color_data = 12'h0ae;
			{8'd46, 8'd5}: color_data = 12'h09d;
			{8'd46, 8'd6}: color_data = 12'h09d;
			{8'd46, 8'd7}: color_data = 12'h09d;
			{8'd46, 8'd8}: color_data = 12'h09d;
			{8'd46, 8'd9}: color_data = 12'h09d;
			{8'd46, 8'd10}: color_data = 12'h0ae;
			{8'd46, 8'd11}: color_data = 12'h069;
			{8'd46, 8'd12}: color_data = 12'h000;
			{8'd46, 8'd13}: color_data = 12'h000;
			{8'd46, 8'd14}: color_data = 12'h000;
			{8'd46, 8'd15}: color_data = 12'h000;
			{8'd46, 8'd16}: color_data = 12'h069;
			{8'd46, 8'd17}: color_data = 12'h0ae;
			{8'd46, 8'd18}: color_data = 12'h09d;
			{8'd46, 8'd19}: color_data = 12'h09d;
			{8'd46, 8'd20}: color_data = 12'h09d;
			{8'd46, 8'd21}: color_data = 12'h09d;
			{8'd46, 8'd22}: color_data = 12'h09d;
			{8'd46, 8'd23}: color_data = 12'h09d;
			{8'd46, 8'd24}: color_data = 12'h09d;
			{8'd46, 8'd25}: color_data = 12'h09d;
			{8'd46, 8'd26}: color_data = 12'h09d;
			{8'd46, 8'd27}: color_data = 12'h09d;
			{8'd46, 8'd28}: color_data = 12'h09d;
			{8'd46, 8'd29}: color_data = 12'h08c;
			{8'd46, 8'd30}: color_data = 12'h000;
			{8'd46, 8'd31}: color_data = 12'h000;
			{8'd46, 8'd32}: color_data = 12'h000;
			{8'd46, 8'd33}: color_data = 12'h000;
			{8'd46, 8'd34}: color_data = 12'h000;
			{8'd46, 8'd35}: color_data = 12'h300;
			{8'd46, 8'd36}: color_data = 12'hb10;
			{8'd46, 8'd37}: color_data = 12'hd20;
			{8'd46, 8'd38}: color_data = 12'he21;
			{8'd46, 8'd39}: color_data = 12'he21;
			{8'd46, 8'd40}: color_data = 12'he21;
			{8'd46, 8'd41}: color_data = 12'he21;
			{8'd46, 8'd42}: color_data = 12'he21;
			{8'd46, 8'd43}: color_data = 12'he21;
			{8'd46, 8'd44}: color_data = 12'he21;
			{8'd46, 8'd45}: color_data = 12'he21;
			{8'd46, 8'd46}: color_data = 12'he21;
			{8'd46, 8'd47}: color_data = 12'he21;
			{8'd46, 8'd48}: color_data = 12'he21;
			{8'd46, 8'd49}: color_data = 12'he21;
			{8'd46, 8'd50}: color_data = 12'he21;
			{8'd46, 8'd51}: color_data = 12'he21;
			{8'd46, 8'd52}: color_data = 12'he21;
			{8'd46, 8'd53}: color_data = 12'he21;
			{8'd46, 8'd54}: color_data = 12'he21;
			{8'd46, 8'd55}: color_data = 12'he21;
			{8'd46, 8'd56}: color_data = 12'he21;
			{8'd46, 8'd57}: color_data = 12'he21;
			{8'd46, 8'd58}: color_data = 12'he21;
			{8'd46, 8'd59}: color_data = 12'he21;
			{8'd46, 8'd60}: color_data = 12'he21;
			{8'd46, 8'd61}: color_data = 12'he21;
			{8'd46, 8'd62}: color_data = 12'he21;
			{8'd46, 8'd63}: color_data = 12'he21;
			{8'd46, 8'd64}: color_data = 12'he21;
			{8'd46, 8'd65}: color_data = 12'he21;
			{8'd46, 8'd66}: color_data = 12'he21;
			{8'd46, 8'd67}: color_data = 12'hb10;
			{8'd46, 8'd68}: color_data = 12'h000;
			{8'd46, 8'd69}: color_data = 12'h000;
			{8'd46, 8'd70}: color_data = 12'h000;
			{8'd46, 8'd71}: color_data = 12'h000;
			{8'd46, 8'd72}: color_data = 12'h000;
			{8'd46, 8'd73}: color_data = 12'h000;
			{8'd46, 8'd74}: color_data = 12'h000;
			{8'd46, 8'd100}: color_data = 12'he00;
			{8'd46, 8'd101}: color_data = 12'hf01;
			{8'd46, 8'd102}: color_data = 12'he00;
			{8'd46, 8'd103}: color_data = 12'he00;
			{8'd46, 8'd104}: color_data = 12'he00;
			{8'd46, 8'd105}: color_data = 12'he00;
			{8'd46, 8'd106}: color_data = 12'hc00;
			{8'd46, 8'd111}: color_data = 12'he00;
			{8'd46, 8'd112}: color_data = 12'he00;
			{8'd46, 8'd113}: color_data = 12'he00;
			{8'd46, 8'd114}: color_data = 12'he01;
			{8'd46, 8'd115}: color_data = 12'he00;
			{8'd46, 8'd116}: color_data = 12'he00;
			{8'd46, 8'd117}: color_data = 12'he00;
			{8'd46, 8'd118}: color_data = 12'he00;
			{8'd46, 8'd119}: color_data = 12'he00;
			{8'd46, 8'd120}: color_data = 12'he00;
			{8'd46, 8'd121}: color_data = 12'he00;
			{8'd46, 8'd122}: color_data = 12'he00;
			{8'd46, 8'd123}: color_data = 12'he00;
			{8'd46, 8'd124}: color_data = 12'he00;
			{8'd46, 8'd125}: color_data = 12'he00;
			{8'd46, 8'd126}: color_data = 12'he01;
			{8'd46, 8'd127}: color_data = 12'he00;
			{8'd46, 8'd128}: color_data = 12'he00;
			{8'd46, 8'd129}: color_data = 12'he00;
			{8'd46, 8'd130}: color_data = 12'he00;
			{8'd46, 8'd131}: color_data = 12'hf00;
			{8'd46, 8'd138}: color_data = 12'he00;
			{8'd46, 8'd139}: color_data = 12'he00;
			{8'd46, 8'd140}: color_data = 12'he00;
			{8'd46, 8'd141}: color_data = 12'he00;
			{8'd46, 8'd142}: color_data = 12'he00;
			{8'd46, 8'd143}: color_data = 12'he01;
			{8'd46, 8'd144}: color_data = 12'he00;
			{8'd47, 8'd1}: color_data = 12'h000;
			{8'd47, 8'd2}: color_data = 12'h000;
			{8'd47, 8'd3}: color_data = 12'h000;
			{8'd47, 8'd4}: color_data = 12'h07a;
			{8'd47, 8'd5}: color_data = 12'h0ae;
			{8'd47, 8'd6}: color_data = 12'h09d;
			{8'd47, 8'd7}: color_data = 12'h09d;
			{8'd47, 8'd8}: color_data = 12'h09d;
			{8'd47, 8'd9}: color_data = 12'h09d;
			{8'd47, 8'd10}: color_data = 12'h09d;
			{8'd47, 8'd11}: color_data = 12'h0ae;
			{8'd47, 8'd12}: color_data = 12'h045;
			{8'd47, 8'd13}: color_data = 12'h000;
			{8'd47, 8'd14}: color_data = 12'h000;
			{8'd47, 8'd15}: color_data = 12'h000;
			{8'd47, 8'd16}: color_data = 12'h011;
			{8'd47, 8'd17}: color_data = 12'h08c;
			{8'd47, 8'd18}: color_data = 12'h09d;
			{8'd47, 8'd19}: color_data = 12'h09d;
			{8'd47, 8'd20}: color_data = 12'h09d;
			{8'd47, 8'd21}: color_data = 12'h09d;
			{8'd47, 8'd22}: color_data = 12'h09d;
			{8'd47, 8'd23}: color_data = 12'h09d;
			{8'd47, 8'd24}: color_data = 12'h09d;
			{8'd47, 8'd25}: color_data = 12'h09d;
			{8'd47, 8'd26}: color_data = 12'h09d;
			{8'd47, 8'd27}: color_data = 12'h0ae;
			{8'd47, 8'd28}: color_data = 12'h0ae;
			{8'd47, 8'd29}: color_data = 12'h069;
			{8'd47, 8'd30}: color_data = 12'h000;
			{8'd47, 8'd31}: color_data = 12'h000;
			{8'd47, 8'd32}: color_data = 12'h000;
			{8'd47, 8'd33}: color_data = 12'h000;
			{8'd47, 8'd34}: color_data = 12'h000;
			{8'd47, 8'd35}: color_data = 12'h000;
			{8'd47, 8'd36}: color_data = 12'h000;
			{8'd47, 8'd37}: color_data = 12'h100;
			{8'd47, 8'd38}: color_data = 12'h300;
			{8'd47, 8'd39}: color_data = 12'h600;
			{8'd47, 8'd40}: color_data = 12'h910;
			{8'd47, 8'd41}: color_data = 12'hb10;
			{8'd47, 8'd42}: color_data = 12'hd20;
			{8'd47, 8'd43}: color_data = 12'he21;
			{8'd47, 8'd44}: color_data = 12'he21;
			{8'd47, 8'd45}: color_data = 12'he21;
			{8'd47, 8'd46}: color_data = 12'he21;
			{8'd47, 8'd47}: color_data = 12'he21;
			{8'd47, 8'd48}: color_data = 12'he21;
			{8'd47, 8'd49}: color_data = 12'he21;
			{8'd47, 8'd50}: color_data = 12'he21;
			{8'd47, 8'd51}: color_data = 12'he21;
			{8'd47, 8'd52}: color_data = 12'he21;
			{8'd47, 8'd53}: color_data = 12'he21;
			{8'd47, 8'd54}: color_data = 12'he21;
			{8'd47, 8'd55}: color_data = 12'he21;
			{8'd47, 8'd56}: color_data = 12'he21;
			{8'd47, 8'd57}: color_data = 12'he21;
			{8'd47, 8'd58}: color_data = 12'he21;
			{8'd47, 8'd59}: color_data = 12'he21;
			{8'd47, 8'd60}: color_data = 12'he21;
			{8'd47, 8'd61}: color_data = 12'he21;
			{8'd47, 8'd62}: color_data = 12'he21;
			{8'd47, 8'd63}: color_data = 12'he21;
			{8'd47, 8'd64}: color_data = 12'he21;
			{8'd47, 8'd65}: color_data = 12'he21;
			{8'd47, 8'd66}: color_data = 12'he21;
			{8'd47, 8'd67}: color_data = 12'h910;
			{8'd47, 8'd68}: color_data = 12'h000;
			{8'd47, 8'd69}: color_data = 12'h000;
			{8'd47, 8'd70}: color_data = 12'h000;
			{8'd47, 8'd71}: color_data = 12'h000;
			{8'd47, 8'd72}: color_data = 12'h000;
			{8'd47, 8'd73}: color_data = 12'h000;
			{8'd47, 8'd74}: color_data = 12'h000;
			{8'd47, 8'd100}: color_data = 12'he00;
			{8'd47, 8'd101}: color_data = 12'hf01;
			{8'd47, 8'd102}: color_data = 12'he00;
			{8'd47, 8'd103}: color_data = 12'he00;
			{8'd47, 8'd104}: color_data = 12'he00;
			{8'd47, 8'd105}: color_data = 12'he00;
			{8'd47, 8'd106}: color_data = 12'hc00;
			{8'd47, 8'd111}: color_data = 12'he01;
			{8'd47, 8'd112}: color_data = 12'he00;
			{8'd47, 8'd113}: color_data = 12'he00;
			{8'd47, 8'd114}: color_data = 12'he00;
			{8'd47, 8'd115}: color_data = 12'he00;
			{8'd47, 8'd116}: color_data = 12'he00;
			{8'd47, 8'd117}: color_data = 12'he00;
			{8'd47, 8'd118}: color_data = 12'he00;
			{8'd47, 8'd119}: color_data = 12'he00;
			{8'd47, 8'd120}: color_data = 12'he00;
			{8'd47, 8'd121}: color_data = 12'he00;
			{8'd47, 8'd122}: color_data = 12'he00;
			{8'd47, 8'd123}: color_data = 12'he00;
			{8'd47, 8'd124}: color_data = 12'he00;
			{8'd47, 8'd125}: color_data = 12'he00;
			{8'd47, 8'd126}: color_data = 12'he00;
			{8'd47, 8'd127}: color_data = 12'he01;
			{8'd47, 8'd128}: color_data = 12'hd00;
			{8'd47, 8'd138}: color_data = 12'he00;
			{8'd47, 8'd139}: color_data = 12'he00;
			{8'd47, 8'd140}: color_data = 12'he00;
			{8'd47, 8'd141}: color_data = 12'he00;
			{8'd47, 8'd142}: color_data = 12'he00;
			{8'd47, 8'd143}: color_data = 12'he01;
			{8'd47, 8'd144}: color_data = 12'he00;
			{8'd48, 8'd1}: color_data = 12'h000;
			{8'd48, 8'd2}: color_data = 12'h000;
			{8'd48, 8'd3}: color_data = 12'h000;
			{8'd48, 8'd4}: color_data = 12'h012;
			{8'd48, 8'd5}: color_data = 12'h08c;
			{8'd48, 8'd6}: color_data = 12'h09d;
			{8'd48, 8'd7}: color_data = 12'h09d;
			{8'd48, 8'd8}: color_data = 12'h09d;
			{8'd48, 8'd9}: color_data = 12'h09d;
			{8'd48, 8'd10}: color_data = 12'h09d;
			{8'd48, 8'd11}: color_data = 12'h09d;
			{8'd48, 8'd12}: color_data = 12'h09d;
			{8'd48, 8'd13}: color_data = 12'h012;
			{8'd48, 8'd14}: color_data = 12'h000;
			{8'd48, 8'd15}: color_data = 12'h000;
			{8'd48, 8'd16}: color_data = 12'h000;
			{8'd48, 8'd17}: color_data = 12'h035;
			{8'd48, 8'd18}: color_data = 12'h09d;
			{8'd48, 8'd19}: color_data = 12'h09d;
			{8'd48, 8'd20}: color_data = 12'h09d;
			{8'd48, 8'd21}: color_data = 12'h09d;
			{8'd48, 8'd22}: color_data = 12'h09d;
			{8'd48, 8'd23}: color_data = 12'h09d;
			{8'd48, 8'd24}: color_data = 12'h09d;
			{8'd48, 8'd25}: color_data = 12'h0ae;
			{8'd48, 8'd26}: color_data = 12'h09d;
			{8'd48, 8'd27}: color_data = 12'h07a;
			{8'd48, 8'd28}: color_data = 12'h034;
			{8'd48, 8'd29}: color_data = 12'h000;
			{8'd48, 8'd30}: color_data = 12'h000;
			{8'd48, 8'd31}: color_data = 12'h000;
			{8'd48, 8'd32}: color_data = 12'h000;
			{8'd48, 8'd33}: color_data = 12'h000;
			{8'd48, 8'd34}: color_data = 12'h000;
			{8'd48, 8'd35}: color_data = 12'h000;
			{8'd48, 8'd36}: color_data = 12'h000;
			{8'd48, 8'd37}: color_data = 12'h000;
			{8'd48, 8'd38}: color_data = 12'h000;
			{8'd48, 8'd39}: color_data = 12'h000;
			{8'd48, 8'd40}: color_data = 12'h000;
			{8'd48, 8'd41}: color_data = 12'h000;
			{8'd48, 8'd42}: color_data = 12'h100;
			{8'd48, 8'd43}: color_data = 12'h300;
			{8'd48, 8'd44}: color_data = 12'h600;
			{8'd48, 8'd45}: color_data = 12'h910;
			{8'd48, 8'd46}: color_data = 12'hb10;
			{8'd48, 8'd47}: color_data = 12'hd20;
			{8'd48, 8'd48}: color_data = 12'he21;
			{8'd48, 8'd49}: color_data = 12'he21;
			{8'd48, 8'd50}: color_data = 12'he21;
			{8'd48, 8'd51}: color_data = 12'he21;
			{8'd48, 8'd52}: color_data = 12'he21;
			{8'd48, 8'd53}: color_data = 12'he21;
			{8'd48, 8'd54}: color_data = 12'he21;
			{8'd48, 8'd55}: color_data = 12'he21;
			{8'd48, 8'd56}: color_data = 12'he21;
			{8'd48, 8'd57}: color_data = 12'he21;
			{8'd48, 8'd58}: color_data = 12'he21;
			{8'd48, 8'd59}: color_data = 12'he21;
			{8'd48, 8'd60}: color_data = 12'he21;
			{8'd48, 8'd61}: color_data = 12'he21;
			{8'd48, 8'd62}: color_data = 12'he21;
			{8'd48, 8'd63}: color_data = 12'he21;
			{8'd48, 8'd64}: color_data = 12'he21;
			{8'd48, 8'd65}: color_data = 12'he21;
			{8'd48, 8'd66}: color_data = 12'he21;
			{8'd48, 8'd67}: color_data = 12'h610;
			{8'd48, 8'd68}: color_data = 12'h000;
			{8'd48, 8'd69}: color_data = 12'h000;
			{8'd48, 8'd70}: color_data = 12'h000;
			{8'd48, 8'd71}: color_data = 12'h000;
			{8'd48, 8'd72}: color_data = 12'h000;
			{8'd48, 8'd73}: color_data = 12'h000;
			{8'd48, 8'd74}: color_data = 12'h000;
			{8'd48, 8'd100}: color_data = 12'he00;
			{8'd48, 8'd101}: color_data = 12'hf01;
			{8'd48, 8'd102}: color_data = 12'he00;
			{8'd48, 8'd103}: color_data = 12'he00;
			{8'd48, 8'd104}: color_data = 12'he00;
			{8'd48, 8'd105}: color_data = 12'he00;
			{8'd48, 8'd106}: color_data = 12'hc00;
			{8'd48, 8'd111}: color_data = 12'he01;
			{8'd48, 8'd112}: color_data = 12'he00;
			{8'd48, 8'd113}: color_data = 12'he00;
			{8'd48, 8'd114}: color_data = 12'he00;
			{8'd48, 8'd115}: color_data = 12'he00;
			{8'd48, 8'd116}: color_data = 12'he00;
			{8'd48, 8'd117}: color_data = 12'he00;
			{8'd48, 8'd118}: color_data = 12'he00;
			{8'd48, 8'd119}: color_data = 12'he00;
			{8'd48, 8'd120}: color_data = 12'he00;
			{8'd48, 8'd121}: color_data = 12'he01;
			{8'd48, 8'd122}: color_data = 12'he00;
			{8'd48, 8'd123}: color_data = 12'he00;
			{8'd48, 8'd124}: color_data = 12'he00;
			{8'd48, 8'd125}: color_data = 12'hd00;
			{8'd48, 8'd138}: color_data = 12'he00;
			{8'd48, 8'd139}: color_data = 12'he00;
			{8'd48, 8'd140}: color_data = 12'he00;
			{8'd48, 8'd141}: color_data = 12'he00;
			{8'd48, 8'd142}: color_data = 12'he00;
			{8'd48, 8'd143}: color_data = 12'he01;
			{8'd48, 8'd144}: color_data = 12'he00;
			{8'd49, 8'd2}: color_data = 12'h000;
			{8'd49, 8'd3}: color_data = 12'h000;
			{8'd49, 8'd4}: color_data = 12'h000;
			{8'd49, 8'd5}: color_data = 12'h034;
			{8'd49, 8'd6}: color_data = 12'h09d;
			{8'd49, 8'd7}: color_data = 12'h09d;
			{8'd49, 8'd8}: color_data = 12'h09d;
			{8'd49, 8'd9}: color_data = 12'h09d;
			{8'd49, 8'd10}: color_data = 12'h09d;
			{8'd49, 8'd11}: color_data = 12'h0ae;
			{8'd49, 8'd12}: color_data = 12'h069;
			{8'd49, 8'd13}: color_data = 12'h001;
			{8'd49, 8'd14}: color_data = 12'h000;
			{8'd49, 8'd15}: color_data = 12'h000;
			{8'd49, 8'd16}: color_data = 12'h000;
			{8'd49, 8'd17}: color_data = 12'h000;
			{8'd49, 8'd18}: color_data = 12'h069;
			{8'd49, 8'd19}: color_data = 12'h0ae;
			{8'd49, 8'd20}: color_data = 12'h09d;
			{8'd49, 8'd21}: color_data = 12'h09d;
			{8'd49, 8'd22}: color_data = 12'h09d;
			{8'd49, 8'd23}: color_data = 12'h0ae;
			{8'd49, 8'd24}: color_data = 12'h09d;
			{8'd49, 8'd25}: color_data = 12'h068;
			{8'd49, 8'd26}: color_data = 12'h023;
			{8'd49, 8'd27}: color_data = 12'h000;
			{8'd49, 8'd28}: color_data = 12'h000;
			{8'd49, 8'd29}: color_data = 12'h000;
			{8'd49, 8'd30}: color_data = 12'h000;
			{8'd49, 8'd31}: color_data = 12'h000;
			{8'd49, 8'd32}: color_data = 12'h000;
			{8'd49, 8'd33}: color_data = 12'h000;
			{8'd49, 8'd34}: color_data = 12'h000;
			{8'd49, 8'd35}: color_data = 12'h000;
			{8'd49, 8'd36}: color_data = 12'h000;
			{8'd49, 8'd37}: color_data = 12'h000;
			{8'd49, 8'd38}: color_data = 12'h000;
			{8'd49, 8'd39}: color_data = 12'h000;
			{8'd49, 8'd40}: color_data = 12'h000;
			{8'd49, 8'd41}: color_data = 12'h000;
			{8'd49, 8'd42}: color_data = 12'h000;
			{8'd49, 8'd43}: color_data = 12'h000;
			{8'd49, 8'd44}: color_data = 12'h000;
			{8'd49, 8'd45}: color_data = 12'h000;
			{8'd49, 8'd46}: color_data = 12'h000;
			{8'd49, 8'd47}: color_data = 12'h100;
			{8'd49, 8'd48}: color_data = 12'h300;
			{8'd49, 8'd49}: color_data = 12'h610;
			{8'd49, 8'd50}: color_data = 12'h910;
			{8'd49, 8'd51}: color_data = 12'hb10;
			{8'd49, 8'd52}: color_data = 12'hd20;
			{8'd49, 8'd53}: color_data = 12'he21;
			{8'd49, 8'd54}: color_data = 12'he21;
			{8'd49, 8'd55}: color_data = 12'he21;
			{8'd49, 8'd56}: color_data = 12'he21;
			{8'd49, 8'd57}: color_data = 12'he21;
			{8'd49, 8'd58}: color_data = 12'he21;
			{8'd49, 8'd59}: color_data = 12'he21;
			{8'd49, 8'd60}: color_data = 12'he21;
			{8'd49, 8'd61}: color_data = 12'he21;
			{8'd49, 8'd62}: color_data = 12'he21;
			{8'd49, 8'd63}: color_data = 12'he21;
			{8'd49, 8'd64}: color_data = 12'he21;
			{8'd49, 8'd65}: color_data = 12'he21;
			{8'd49, 8'd66}: color_data = 12'he21;
			{8'd49, 8'd67}: color_data = 12'h300;
			{8'd49, 8'd68}: color_data = 12'h000;
			{8'd49, 8'd69}: color_data = 12'h000;
			{8'd49, 8'd70}: color_data = 12'h000;
			{8'd49, 8'd71}: color_data = 12'h000;
			{8'd49, 8'd72}: color_data = 12'h000;
			{8'd49, 8'd73}: color_data = 12'h000;
			{8'd49, 8'd74}: color_data = 12'h000;
			{8'd49, 8'd100}: color_data = 12'he00;
			{8'd49, 8'd101}: color_data = 12'hf01;
			{8'd49, 8'd102}: color_data = 12'he00;
			{8'd49, 8'd103}: color_data = 12'he00;
			{8'd49, 8'd104}: color_data = 12'he00;
			{8'd49, 8'd105}: color_data = 12'he00;
			{8'd49, 8'd106}: color_data = 12'hc00;
			{8'd49, 8'd111}: color_data = 12'he00;
			{8'd49, 8'd112}: color_data = 12'he00;
			{8'd49, 8'd113}: color_data = 12'he00;
			{8'd49, 8'd114}: color_data = 12'he00;
			{8'd49, 8'd115}: color_data = 12'he00;
			{8'd49, 8'd116}: color_data = 12'he00;
			{8'd49, 8'd117}: color_data = 12'he00;
			{8'd49, 8'd118}: color_data = 12'he01;
			{8'd49, 8'd119}: color_data = 12'he00;
			{8'd49, 8'd120}: color_data = 12'he00;
			{8'd49, 8'd121}: color_data = 12'he00;
			{8'd49, 8'd122}: color_data = 12'he00;
			{8'd49, 8'd138}: color_data = 12'he00;
			{8'd49, 8'd139}: color_data = 12'he00;
			{8'd49, 8'd140}: color_data = 12'he00;
			{8'd49, 8'd141}: color_data = 12'he00;
			{8'd49, 8'd142}: color_data = 12'he00;
			{8'd49, 8'd143}: color_data = 12'he01;
			{8'd49, 8'd144}: color_data = 12'he00;
			{8'd50, 8'd3}: color_data = 12'h000;
			{8'd50, 8'd4}: color_data = 12'h000;
			{8'd50, 8'd5}: color_data = 12'h000;
			{8'd50, 8'd6}: color_data = 12'h046;
			{8'd50, 8'd7}: color_data = 12'h0ae;
			{8'd50, 8'd8}: color_data = 12'h09d;
			{8'd50, 8'd9}: color_data = 12'h09d;
			{8'd50, 8'd10}: color_data = 12'h09d;
			{8'd50, 8'd11}: color_data = 12'h057;
			{8'd50, 8'd12}: color_data = 12'h000;
			{8'd50, 8'd13}: color_data = 12'h000;
			{8'd50, 8'd14}: color_data = 12'h000;
			{8'd50, 8'd15}: color_data = 12'h000;
			{8'd50, 8'd16}: color_data = 12'h000;
			{8'd50, 8'd17}: color_data = 12'h000;
			{8'd50, 8'd18}: color_data = 12'h012;
			{8'd50, 8'd19}: color_data = 12'h09c;
			{8'd50, 8'd20}: color_data = 12'h0ae;
			{8'd50, 8'd21}: color_data = 12'h0ae;
			{8'd50, 8'd22}: color_data = 12'h08c;
			{8'd50, 8'd23}: color_data = 12'h057;
			{8'd50, 8'd24}: color_data = 12'h011;
			{8'd50, 8'd25}: color_data = 12'h000;
			{8'd50, 8'd26}: color_data = 12'h000;
			{8'd50, 8'd27}: color_data = 12'h000;
			{8'd50, 8'd28}: color_data = 12'h000;
			{8'd50, 8'd29}: color_data = 12'h000;
			{8'd50, 8'd30}: color_data = 12'h000;
			{8'd50, 8'd31}: color_data = 12'h000;
			{8'd50, 8'd32}: color_data = 12'h000;
			{8'd50, 8'd33}: color_data = 12'h000;
			{8'd50, 8'd34}: color_data = 12'h000;
			{8'd50, 8'd35}: color_data = 12'h000;
			{8'd50, 8'd36}: color_data = 12'h000;
			{8'd50, 8'd37}: color_data = 12'h000;
			{8'd50, 8'd38}: color_data = 12'h000;
			{8'd50, 8'd39}: color_data = 12'h000;
			{8'd50, 8'd40}: color_data = 12'h000;
			{8'd50, 8'd41}: color_data = 12'h000;
			{8'd50, 8'd42}: color_data = 12'h000;
			{8'd50, 8'd43}: color_data = 12'h000;
			{8'd50, 8'd44}: color_data = 12'h000;
			{8'd50, 8'd45}: color_data = 12'h000;
			{8'd50, 8'd46}: color_data = 12'h000;
			{8'd50, 8'd47}: color_data = 12'h000;
			{8'd50, 8'd48}: color_data = 12'h000;
			{8'd50, 8'd49}: color_data = 12'h000;
			{8'd50, 8'd50}: color_data = 12'h000;
			{8'd50, 8'd51}: color_data = 12'h000;
			{8'd50, 8'd52}: color_data = 12'h100;
			{8'd50, 8'd53}: color_data = 12'h300;
			{8'd50, 8'd54}: color_data = 12'h610;
			{8'd50, 8'd55}: color_data = 12'h910;
			{8'd50, 8'd56}: color_data = 12'hb10;
			{8'd50, 8'd57}: color_data = 12'hd20;
			{8'd50, 8'd58}: color_data = 12'he21;
			{8'd50, 8'd59}: color_data = 12'he21;
			{8'd50, 8'd60}: color_data = 12'he21;
			{8'd50, 8'd61}: color_data = 12'he21;
			{8'd50, 8'd62}: color_data = 12'he21;
			{8'd50, 8'd63}: color_data = 12'he21;
			{8'd50, 8'd64}: color_data = 12'he21;
			{8'd50, 8'd65}: color_data = 12'he21;
			{8'd50, 8'd66}: color_data = 12'hd20;
			{8'd50, 8'd67}: color_data = 12'h100;
			{8'd50, 8'd68}: color_data = 12'h000;
			{8'd50, 8'd69}: color_data = 12'h000;
			{8'd50, 8'd70}: color_data = 12'h000;
			{8'd50, 8'd71}: color_data = 12'h000;
			{8'd50, 8'd72}: color_data = 12'h000;
			{8'd50, 8'd73}: color_data = 12'h000;
			{8'd50, 8'd74}: color_data = 12'h000;
			{8'd50, 8'd100}: color_data = 12'he00;
			{8'd50, 8'd101}: color_data = 12'hf01;
			{8'd50, 8'd102}: color_data = 12'he00;
			{8'd50, 8'd103}: color_data = 12'he00;
			{8'd50, 8'd104}: color_data = 12'he00;
			{8'd50, 8'd105}: color_data = 12'he00;
			{8'd50, 8'd106}: color_data = 12'hc00;
			{8'd50, 8'd111}: color_data = 12'he00;
			{8'd50, 8'd112}: color_data = 12'he00;
			{8'd50, 8'd113}: color_data = 12'he00;
			{8'd50, 8'd114}: color_data = 12'he00;
			{8'd50, 8'd115}: color_data = 12'he00;
			{8'd50, 8'd116}: color_data = 12'he00;
			{8'd50, 8'd117}: color_data = 12'he00;
			{8'd50, 8'd118}: color_data = 12'he00;
			{8'd50, 8'd119}: color_data = 12'he01;
			{8'd50, 8'd120}: color_data = 12'hc00;
			{8'd50, 8'd138}: color_data = 12'he00;
			{8'd50, 8'd139}: color_data = 12'he00;
			{8'd50, 8'd140}: color_data = 12'he00;
			{8'd50, 8'd141}: color_data = 12'he00;
			{8'd50, 8'd142}: color_data = 12'he00;
			{8'd50, 8'd143}: color_data = 12'he01;
			{8'd50, 8'd144}: color_data = 12'he00;
			{8'd51, 8'd3}: color_data = 12'h000;
			{8'd51, 8'd4}: color_data = 12'h000;
			{8'd51, 8'd5}: color_data = 12'h000;
			{8'd51, 8'd6}: color_data = 12'h000;
			{8'd51, 8'd7}: color_data = 12'h069;
			{8'd51, 8'd8}: color_data = 12'h0ae;
			{8'd51, 8'd9}: color_data = 12'h09c;
			{8'd51, 8'd10}: color_data = 12'h034;
			{8'd51, 8'd11}: color_data = 12'h000;
			{8'd51, 8'd12}: color_data = 12'h000;
			{8'd51, 8'd13}: color_data = 12'h000;
			{8'd51, 8'd14}: color_data = 12'h000;
			{8'd51, 8'd15}: color_data = 12'h000;
			{8'd51, 8'd16}: color_data = 12'h000;
			{8'd51, 8'd17}: color_data = 12'h000;
			{8'd51, 8'd18}: color_data = 12'h000;
			{8'd51, 8'd19}: color_data = 12'h035;
			{8'd51, 8'd20}: color_data = 12'h08b;
			{8'd51, 8'd21}: color_data = 12'h045;
			{8'd51, 8'd22}: color_data = 12'h001;
			{8'd51, 8'd23}: color_data = 12'h000;
			{8'd51, 8'd24}: color_data = 12'h000;
			{8'd51, 8'd25}: color_data = 12'h000;
			{8'd51, 8'd26}: color_data = 12'h000;
			{8'd51, 8'd27}: color_data = 12'h000;
			{8'd51, 8'd28}: color_data = 12'h000;
			{8'd51, 8'd29}: color_data = 12'h000;
			{8'd51, 8'd30}: color_data = 12'h000;
			{8'd51, 8'd31}: color_data = 12'h000;
			{8'd51, 8'd32}: color_data = 12'h000;
			{8'd51, 8'd33}: color_data = 12'h000;
			{8'd51, 8'd34}: color_data = 12'h000;
			{8'd51, 8'd35}: color_data = 12'h000;
			{8'd51, 8'd36}: color_data = 12'h000;
			{8'd51, 8'd37}: color_data = 12'h000;
			{8'd51, 8'd38}: color_data = 12'h000;
			{8'd51, 8'd39}: color_data = 12'h000;
			{8'd51, 8'd40}: color_data = 12'h000;
			{8'd51, 8'd41}: color_data = 12'h000;
			{8'd51, 8'd42}: color_data = 12'h000;
			{8'd51, 8'd43}: color_data = 12'h000;
			{8'd51, 8'd44}: color_data = 12'h000;
			{8'd51, 8'd45}: color_data = 12'h000;
			{8'd51, 8'd46}: color_data = 12'h000;
			{8'd51, 8'd47}: color_data = 12'h000;
			{8'd51, 8'd48}: color_data = 12'h000;
			{8'd51, 8'd49}: color_data = 12'h000;
			{8'd51, 8'd50}: color_data = 12'h000;
			{8'd51, 8'd51}: color_data = 12'h000;
			{8'd51, 8'd52}: color_data = 12'h000;
			{8'd51, 8'd53}: color_data = 12'h000;
			{8'd51, 8'd54}: color_data = 12'h000;
			{8'd51, 8'd55}: color_data = 12'h000;
			{8'd51, 8'd56}: color_data = 12'h000;
			{8'd51, 8'd57}: color_data = 12'h100;
			{8'd51, 8'd58}: color_data = 12'h400;
			{8'd51, 8'd59}: color_data = 12'h610;
			{8'd51, 8'd60}: color_data = 12'h910;
			{8'd51, 8'd61}: color_data = 12'hc10;
			{8'd51, 8'd62}: color_data = 12'hd20;
			{8'd51, 8'd63}: color_data = 12'he21;
			{8'd51, 8'd64}: color_data = 12'he21;
			{8'd51, 8'd65}: color_data = 12'hf21;
			{8'd51, 8'd66}: color_data = 12'hb10;
			{8'd51, 8'd67}: color_data = 12'h000;
			{8'd51, 8'd68}: color_data = 12'h000;
			{8'd51, 8'd69}: color_data = 12'h000;
			{8'd51, 8'd70}: color_data = 12'h000;
			{8'd51, 8'd71}: color_data = 12'h000;
			{8'd51, 8'd72}: color_data = 12'h000;
			{8'd51, 8'd73}: color_data = 12'h000;
			{8'd51, 8'd100}: color_data = 12'he00;
			{8'd51, 8'd101}: color_data = 12'hf01;
			{8'd51, 8'd102}: color_data = 12'he00;
			{8'd51, 8'd103}: color_data = 12'he00;
			{8'd51, 8'd104}: color_data = 12'he00;
			{8'd51, 8'd105}: color_data = 12'he00;
			{8'd51, 8'd106}: color_data = 12'hc00;
			{8'd51, 8'd111}: color_data = 12'he00;
			{8'd51, 8'd112}: color_data = 12'he00;
			{8'd51, 8'd113}: color_data = 12'hf01;
			{8'd51, 8'd114}: color_data = 12'he00;
			{8'd51, 8'd115}: color_data = 12'he00;
			{8'd51, 8'd116}: color_data = 12'he00;
			{8'd51, 8'd117}: color_data = 12'hd00;
			{8'd51, 8'd138}: color_data = 12'he00;
			{8'd51, 8'd139}: color_data = 12'he00;
			{8'd51, 8'd140}: color_data = 12'he00;
			{8'd51, 8'd141}: color_data = 12'he00;
			{8'd51, 8'd142}: color_data = 12'he00;
			{8'd51, 8'd143}: color_data = 12'he01;
			{8'd51, 8'd144}: color_data = 12'he00;
			{8'd52, 8'd2}: color_data = 12'h000;
			{8'd52, 8'd3}: color_data = 12'h000;
			{8'd52, 8'd4}: color_data = 12'h000;
			{8'd52, 8'd5}: color_data = 12'h000;
			{8'd52, 8'd6}: color_data = 12'h000;
			{8'd52, 8'd7}: color_data = 12'h011;
			{8'd52, 8'd8}: color_data = 12'h069;
			{8'd52, 8'd9}: color_data = 12'h022;
			{8'd52, 8'd10}: color_data = 12'h000;
			{8'd52, 8'd11}: color_data = 12'h000;
			{8'd52, 8'd12}: color_data = 12'h000;
			{8'd52, 8'd13}: color_data = 12'h000;
			{8'd52, 8'd14}: color_data = 12'h000;
			{8'd52, 8'd15}: color_data = 12'h000;
			{8'd52, 8'd16}: color_data = 12'h000;
			{8'd52, 8'd17}: color_data = 12'h000;
			{8'd52, 8'd18}: color_data = 12'h000;
			{8'd52, 8'd19}: color_data = 12'h000;
			{8'd52, 8'd20}: color_data = 12'h000;
			{8'd52, 8'd21}: color_data = 12'h000;
			{8'd52, 8'd22}: color_data = 12'h000;
			{8'd52, 8'd23}: color_data = 12'h110;
			{8'd52, 8'd24}: color_data = 12'h220;
			{8'd52, 8'd25}: color_data = 12'h000;
			{8'd52, 8'd26}: color_data = 12'h000;
			{8'd52, 8'd27}: color_data = 12'h000;
			{8'd52, 8'd28}: color_data = 12'h000;
			{8'd52, 8'd29}: color_data = 12'h000;
			{8'd52, 8'd30}: color_data = 12'h000;
			{8'd52, 8'd31}: color_data = 12'h000;
			{8'd52, 8'd32}: color_data = 12'h000;
			{8'd52, 8'd33}: color_data = 12'h000;
			{8'd52, 8'd34}: color_data = 12'h000;
			{8'd52, 8'd35}: color_data = 12'h000;
			{8'd52, 8'd36}: color_data = 12'h000;
			{8'd52, 8'd37}: color_data = 12'h000;
			{8'd52, 8'd38}: color_data = 12'h000;
			{8'd52, 8'd39}: color_data = 12'h000;
			{8'd52, 8'd40}: color_data = 12'h000;
			{8'd52, 8'd41}: color_data = 12'h000;
			{8'd52, 8'd42}: color_data = 12'h000;
			{8'd52, 8'd43}: color_data = 12'h000;
			{8'd52, 8'd44}: color_data = 12'h000;
			{8'd52, 8'd45}: color_data = 12'h000;
			{8'd52, 8'd46}: color_data = 12'h000;
			{8'd52, 8'd47}: color_data = 12'h000;
			{8'd52, 8'd48}: color_data = 12'h000;
			{8'd52, 8'd49}: color_data = 12'h120;
			{8'd52, 8'd50}: color_data = 12'h251;
			{8'd52, 8'd51}: color_data = 12'h141;
			{8'd52, 8'd52}: color_data = 12'h120;
			{8'd52, 8'd53}: color_data = 12'h010;
			{8'd52, 8'd54}: color_data = 12'h000;
			{8'd52, 8'd55}: color_data = 12'h000;
			{8'd52, 8'd56}: color_data = 12'h000;
			{8'd52, 8'd57}: color_data = 12'h000;
			{8'd52, 8'd58}: color_data = 12'h000;
			{8'd52, 8'd59}: color_data = 12'h000;
			{8'd52, 8'd60}: color_data = 12'h000;
			{8'd52, 8'd61}: color_data = 12'h000;
			{8'd52, 8'd62}: color_data = 12'h100;
			{8'd52, 8'd63}: color_data = 12'h400;
			{8'd52, 8'd64}: color_data = 12'h710;
			{8'd52, 8'd65}: color_data = 12'ha10;
			{8'd52, 8'd66}: color_data = 12'h610;
			{8'd52, 8'd67}: color_data = 12'h000;
			{8'd52, 8'd68}: color_data = 12'h000;
			{8'd52, 8'd69}: color_data = 12'h000;
			{8'd52, 8'd70}: color_data = 12'h000;
			{8'd52, 8'd71}: color_data = 12'h000;
			{8'd52, 8'd72}: color_data = 12'h000;
			{8'd52, 8'd73}: color_data = 12'h000;
			{8'd52, 8'd74}: color_data = 12'h000;
			{8'd52, 8'd100}: color_data = 12'he00;
			{8'd52, 8'd101}: color_data = 12'hf01;
			{8'd52, 8'd102}: color_data = 12'he00;
			{8'd52, 8'd103}: color_data = 12'he00;
			{8'd52, 8'd104}: color_data = 12'he00;
			{8'd52, 8'd105}: color_data = 12'he00;
			{8'd52, 8'd106}: color_data = 12'hc00;
			{8'd52, 8'd111}: color_data = 12'he01;
			{8'd52, 8'd112}: color_data = 12'he00;
			{8'd52, 8'd113}: color_data = 12'he00;
			{8'd52, 8'd114}: color_data = 12'he00;
			{8'd52, 8'd138}: color_data = 12'he00;
			{8'd52, 8'd139}: color_data = 12'he00;
			{8'd52, 8'd140}: color_data = 12'he00;
			{8'd52, 8'd141}: color_data = 12'he00;
			{8'd52, 8'd142}: color_data = 12'he00;
			{8'd52, 8'd143}: color_data = 12'he01;
			{8'd52, 8'd144}: color_data = 12'he00;
			{8'd53, 8'd2}: color_data = 12'h000;
			{8'd53, 8'd3}: color_data = 12'h000;
			{8'd53, 8'd4}: color_data = 12'h000;
			{8'd53, 8'd5}: color_data = 12'h000;
			{8'd53, 8'd6}: color_data = 12'h000;
			{8'd53, 8'd7}: color_data = 12'h000;
			{8'd53, 8'd8}: color_data = 12'h000;
			{8'd53, 8'd9}: color_data = 12'h000;
			{8'd53, 8'd10}: color_data = 12'h100;
			{8'd53, 8'd11}: color_data = 12'h650;
			{8'd53, 8'd12}: color_data = 12'h760;
			{8'd53, 8'd13}: color_data = 12'h870;
			{8'd53, 8'd14}: color_data = 12'h980;
			{8'd53, 8'd15}: color_data = 12'ha80;
			{8'd53, 8'd16}: color_data = 12'hb90;
			{8'd53, 8'd17}: color_data = 12'hca0;
			{8'd53, 8'd18}: color_data = 12'h430;
			{8'd53, 8'd19}: color_data = 12'h000;
			{8'd53, 8'd20}: color_data = 12'h000;
			{8'd53, 8'd21}: color_data = 12'h220;
			{8'd53, 8'd22}: color_data = 12'h970;
			{8'd53, 8'd23}: color_data = 12'hec0;
			{8'd53, 8'd24}: color_data = 12'hfc0;
			{8'd53, 8'd25}: color_data = 12'h540;
			{8'd53, 8'd26}: color_data = 12'h000;
			{8'd53, 8'd27}: color_data = 12'h000;
			{8'd53, 8'd28}: color_data = 12'h000;
			{8'd53, 8'd29}: color_data = 12'h000;
			{8'd53, 8'd30}: color_data = 12'h000;
			{8'd53, 8'd31}: color_data = 12'h000;
			{8'd53, 8'd32}: color_data = 12'h000;
			{8'd53, 8'd33}: color_data = 12'h000;
			{8'd53, 8'd34}: color_data = 12'h000;
			{8'd53, 8'd35}: color_data = 12'h000;
			{8'd53, 8'd36}: color_data = 12'h000;
			{8'd53, 8'd37}: color_data = 12'h000;
			{8'd53, 8'd38}: color_data = 12'h000;
			{8'd53, 8'd39}: color_data = 12'h000;
			{8'd53, 8'd40}: color_data = 12'h000;
			{8'd53, 8'd41}: color_data = 12'h000;
			{8'd53, 8'd42}: color_data = 12'h000;
			{8'd53, 8'd43}: color_data = 12'h000;
			{8'd53, 8'd44}: color_data = 12'h000;
			{8'd53, 8'd45}: color_data = 12'h010;
			{8'd53, 8'd46}: color_data = 12'h131;
			{8'd53, 8'd47}: color_data = 12'h262;
			{8'd53, 8'd48}: color_data = 12'h392;
			{8'd53, 8'd49}: color_data = 12'h4b3;
			{8'd53, 8'd50}: color_data = 12'h4b3;
			{8'd53, 8'd51}: color_data = 12'h4b3;
			{8'd53, 8'd52}: color_data = 12'h4b3;
			{8'd53, 8'd53}: color_data = 12'h4a3;
			{8'd53, 8'd54}: color_data = 12'h382;
			{8'd53, 8'd55}: color_data = 12'h262;
			{8'd53, 8'd56}: color_data = 12'h141;
			{8'd53, 8'd57}: color_data = 12'h120;
			{8'd53, 8'd58}: color_data = 12'h010;
			{8'd53, 8'd59}: color_data = 12'h000;
			{8'd53, 8'd60}: color_data = 12'h000;
			{8'd53, 8'd61}: color_data = 12'h000;
			{8'd53, 8'd62}: color_data = 12'h000;
			{8'd53, 8'd63}: color_data = 12'h000;
			{8'd53, 8'd64}: color_data = 12'h000;
			{8'd53, 8'd65}: color_data = 12'h000;
			{8'd53, 8'd66}: color_data = 12'h000;
			{8'd53, 8'd67}: color_data = 12'h000;
			{8'd53, 8'd68}: color_data = 12'h000;
			{8'd53, 8'd69}: color_data = 12'h000;
			{8'd53, 8'd70}: color_data = 12'h000;
			{8'd53, 8'd71}: color_data = 12'h000;
			{8'd53, 8'd72}: color_data = 12'h000;
			{8'd53, 8'd73}: color_data = 12'h000;
			{8'd53, 8'd74}: color_data = 12'h000;
			{8'd53, 8'd100}: color_data = 12'he00;
			{8'd53, 8'd101}: color_data = 12'hf01;
			{8'd53, 8'd102}: color_data = 12'he00;
			{8'd53, 8'd103}: color_data = 12'he00;
			{8'd53, 8'd104}: color_data = 12'he00;
			{8'd53, 8'd105}: color_data = 12'he00;
			{8'd53, 8'd106}: color_data = 12'hc00;
			{8'd53, 8'd111}: color_data = 12'hf00;
			{8'd53, 8'd112}: color_data = 12'hf00;
			{8'd53, 8'd138}: color_data = 12'he00;
			{8'd53, 8'd139}: color_data = 12'he00;
			{8'd53, 8'd140}: color_data = 12'he00;
			{8'd53, 8'd141}: color_data = 12'he00;
			{8'd53, 8'd142}: color_data = 12'he00;
			{8'd53, 8'd143}: color_data = 12'he01;
			{8'd53, 8'd144}: color_data = 12'he00;
			{8'd54, 8'd3}: color_data = 12'h000;
			{8'd54, 8'd4}: color_data = 12'h000;
			{8'd54, 8'd5}: color_data = 12'h760;
			{8'd54, 8'd6}: color_data = 12'hb90;
			{8'd54, 8'd7}: color_data = 12'h000;
			{8'd54, 8'd8}: color_data = 12'h000;
			{8'd54, 8'd9}: color_data = 12'h210;
			{8'd54, 8'd10}: color_data = 12'hca0;
			{8'd54, 8'd11}: color_data = 12'hfd0;
			{8'd54, 8'd12}: color_data = 12'hfd0;
			{8'd54, 8'd13}: color_data = 12'hfd0;
			{8'd54, 8'd14}: color_data = 12'hfd0;
			{8'd54, 8'd15}: color_data = 12'hfd0;
			{8'd54, 8'd16}: color_data = 12'hfd0;
			{8'd54, 8'd17}: color_data = 12'hfd0;
			{8'd54, 8'd18}: color_data = 12'hec0;
			{8'd54, 8'd19}: color_data = 12'h980;
			{8'd54, 8'd20}: color_data = 12'ha80;
			{8'd54, 8'd21}: color_data = 12'hfc0;
			{8'd54, 8'd22}: color_data = 12'hfd0;
			{8'd54, 8'd23}: color_data = 12'hfd0;
			{8'd54, 8'd24}: color_data = 12'hfd0;
			{8'd54, 8'd25}: color_data = 12'hfc0;
			{8'd54, 8'd26}: color_data = 12'h430;
			{8'd54, 8'd27}: color_data = 12'h000;
			{8'd54, 8'd28}: color_data = 12'h000;
			{8'd54, 8'd29}: color_data = 12'h000;
			{8'd54, 8'd30}: color_data = 12'h000;
			{8'd54, 8'd31}: color_data = 12'h000;
			{8'd54, 8'd32}: color_data = 12'h000;
			{8'd54, 8'd33}: color_data = 12'h000;
			{8'd54, 8'd34}: color_data = 12'h000;
			{8'd54, 8'd35}: color_data = 12'h000;
			{8'd54, 8'd36}: color_data = 12'h000;
			{8'd54, 8'd37}: color_data = 12'h000;
			{8'd54, 8'd38}: color_data = 12'h000;
			{8'd54, 8'd39}: color_data = 12'h000;
			{8'd54, 8'd40}: color_data = 12'h000;
			{8'd54, 8'd41}: color_data = 12'h000;
			{8'd54, 8'd42}: color_data = 12'h020;
			{8'd54, 8'd43}: color_data = 12'h251;
			{8'd54, 8'd44}: color_data = 12'h382;
			{8'd54, 8'd45}: color_data = 12'h4a3;
			{8'd54, 8'd46}: color_data = 12'h4b3;
			{8'd54, 8'd47}: color_data = 12'h4b3;
			{8'd54, 8'd48}: color_data = 12'h4b3;
			{8'd54, 8'd49}: color_data = 12'h4b3;
			{8'd54, 8'd50}: color_data = 12'h4a3;
			{8'd54, 8'd51}: color_data = 12'h4a3;
			{8'd54, 8'd52}: color_data = 12'h4b3;
			{8'd54, 8'd53}: color_data = 12'h4b3;
			{8'd54, 8'd54}: color_data = 12'h4b3;
			{8'd54, 8'd55}: color_data = 12'h4b3;
			{8'd54, 8'd56}: color_data = 12'h4b3;
			{8'd54, 8'd57}: color_data = 12'h4b3;
			{8'd54, 8'd58}: color_data = 12'h3a3;
			{8'd54, 8'd59}: color_data = 12'h382;
			{8'd54, 8'd60}: color_data = 12'h262;
			{8'd54, 8'd61}: color_data = 12'h141;
			{8'd54, 8'd62}: color_data = 12'h120;
			{8'd54, 8'd63}: color_data = 12'h010;
			{8'd54, 8'd64}: color_data = 12'h000;
			{8'd54, 8'd65}: color_data = 12'h000;
			{8'd54, 8'd66}: color_data = 12'h000;
			{8'd54, 8'd67}: color_data = 12'h000;
			{8'd54, 8'd68}: color_data = 12'h000;
			{8'd54, 8'd69}: color_data = 12'h000;
			{8'd54, 8'd70}: color_data = 12'h000;
			{8'd54, 8'd71}: color_data = 12'h000;
			{8'd54, 8'd72}: color_data = 12'h000;
			{8'd54, 8'd73}: color_data = 12'h000;
			{8'd54, 8'd74}: color_data = 12'h000;
			{8'd54, 8'd100}: color_data = 12'he00;
			{8'd54, 8'd101}: color_data = 12'hf01;
			{8'd54, 8'd102}: color_data = 12'he00;
			{8'd54, 8'd103}: color_data = 12'he00;
			{8'd54, 8'd104}: color_data = 12'he00;
			{8'd54, 8'd105}: color_data = 12'he00;
			{8'd54, 8'd106}: color_data = 12'hc00;
			{8'd54, 8'd138}: color_data = 12'he00;
			{8'd54, 8'd139}: color_data = 12'he00;
			{8'd54, 8'd140}: color_data = 12'he00;
			{8'd54, 8'd141}: color_data = 12'he00;
			{8'd54, 8'd142}: color_data = 12'he00;
			{8'd54, 8'd143}: color_data = 12'he01;
			{8'd54, 8'd144}: color_data = 12'he00;
			{8'd55, 8'd3}: color_data = 12'h000;
			{8'd55, 8'd4}: color_data = 12'h000;
			{8'd55, 8'd5}: color_data = 12'h650;
			{8'd55, 8'd6}: color_data = 12'hfd0;
			{8'd55, 8'd7}: color_data = 12'hb90;
			{8'd55, 8'd8}: color_data = 12'h970;
			{8'd55, 8'd9}: color_data = 12'heb0;
			{8'd55, 8'd10}: color_data = 12'hfd0;
			{8'd55, 8'd11}: color_data = 12'hfc0;
			{8'd55, 8'd12}: color_data = 12'hfc0;
			{8'd55, 8'd13}: color_data = 12'hfc0;
			{8'd55, 8'd14}: color_data = 12'hfc0;
			{8'd55, 8'd15}: color_data = 12'hfc0;
			{8'd55, 8'd16}: color_data = 12'hfc0;
			{8'd55, 8'd17}: color_data = 12'hfc0;
			{8'd55, 8'd18}: color_data = 12'hfd0;
			{8'd55, 8'd19}: color_data = 12'hfd0;
			{8'd55, 8'd20}: color_data = 12'hfd0;
			{8'd55, 8'd21}: color_data = 12'hfd0;
			{8'd55, 8'd22}: color_data = 12'hfc0;
			{8'd55, 8'd23}: color_data = 12'hfc0;
			{8'd55, 8'd24}: color_data = 12'hfc0;
			{8'd55, 8'd25}: color_data = 12'hfd0;
			{8'd55, 8'd26}: color_data = 12'hec0;
			{8'd55, 8'd27}: color_data = 12'h320;
			{8'd55, 8'd28}: color_data = 12'h000;
			{8'd55, 8'd29}: color_data = 12'h000;
			{8'd55, 8'd30}: color_data = 12'h000;
			{8'd55, 8'd31}: color_data = 12'h000;
			{8'd55, 8'd32}: color_data = 12'h000;
			{8'd55, 8'd33}: color_data = 12'h000;
			{8'd55, 8'd34}: color_data = 12'h000;
			{8'd55, 8'd35}: color_data = 12'h000;
			{8'd55, 8'd36}: color_data = 12'h000;
			{8'd55, 8'd37}: color_data = 12'h000;
			{8'd55, 8'd38}: color_data = 12'h010;
			{8'd55, 8'd39}: color_data = 12'h131;
			{8'd55, 8'd40}: color_data = 12'h262;
			{8'd55, 8'd41}: color_data = 12'h392;
			{8'd55, 8'd42}: color_data = 12'h4a3;
			{8'd55, 8'd43}: color_data = 12'h4b3;
			{8'd55, 8'd44}: color_data = 12'h4b3;
			{8'd55, 8'd45}: color_data = 12'h4b3;
			{8'd55, 8'd46}: color_data = 12'h4a3;
			{8'd55, 8'd47}: color_data = 12'h4a3;
			{8'd55, 8'd48}: color_data = 12'h4a3;
			{8'd55, 8'd49}: color_data = 12'h4a3;
			{8'd55, 8'd50}: color_data = 12'h4a3;
			{8'd55, 8'd51}: color_data = 12'h4a3;
			{8'd55, 8'd52}: color_data = 12'h4a3;
			{8'd55, 8'd53}: color_data = 12'h4a3;
			{8'd55, 8'd54}: color_data = 12'h4a3;
			{8'd55, 8'd55}: color_data = 12'h4a3;
			{8'd55, 8'd56}: color_data = 12'h4a3;
			{8'd55, 8'd57}: color_data = 12'h4b3;
			{8'd55, 8'd58}: color_data = 12'h4b3;
			{8'd55, 8'd59}: color_data = 12'h4b3;
			{8'd55, 8'd60}: color_data = 12'h4b3;
			{8'd55, 8'd61}: color_data = 12'h4b3;
			{8'd55, 8'd62}: color_data = 12'h4b3;
			{8'd55, 8'd63}: color_data = 12'h3a3;
			{8'd55, 8'd64}: color_data = 12'h382;
			{8'd55, 8'd65}: color_data = 12'h262;
			{8'd55, 8'd66}: color_data = 12'h141;
			{8'd55, 8'd67}: color_data = 12'h010;
			{8'd55, 8'd68}: color_data = 12'h000;
			{8'd55, 8'd69}: color_data = 12'h000;
			{8'd55, 8'd70}: color_data = 12'h000;
			{8'd55, 8'd71}: color_data = 12'h000;
			{8'd55, 8'd72}: color_data = 12'h000;
			{8'd55, 8'd73}: color_data = 12'h000;
			{8'd55, 8'd74}: color_data = 12'h000;
			{8'd55, 8'd100}: color_data = 12'he00;
			{8'd55, 8'd101}: color_data = 12'hf01;
			{8'd55, 8'd102}: color_data = 12'he00;
			{8'd55, 8'd103}: color_data = 12'he00;
			{8'd55, 8'd104}: color_data = 12'he00;
			{8'd55, 8'd105}: color_data = 12'he00;
			{8'd55, 8'd106}: color_data = 12'hc00;
			{8'd55, 8'd111}: color_data = 12'he00;
			{8'd55, 8'd112}: color_data = 12'he00;
			{8'd55, 8'd113}: color_data = 12'he00;
			{8'd55, 8'd114}: color_data = 12'he00;
			{8'd55, 8'd115}: color_data = 12'he00;
			{8'd55, 8'd116}: color_data = 12'hf00;
			{8'd55, 8'd117}: color_data = 12'he00;
			{8'd55, 8'd118}: color_data = 12'he00;
			{8'd55, 8'd119}: color_data = 12'he00;
			{8'd55, 8'd120}: color_data = 12'he00;
			{8'd55, 8'd121}: color_data = 12'he00;
			{8'd55, 8'd122}: color_data = 12'he00;
			{8'd55, 8'd123}: color_data = 12'he00;
			{8'd55, 8'd124}: color_data = 12'he00;
			{8'd55, 8'd125}: color_data = 12'he00;
			{8'd55, 8'd126}: color_data = 12'he00;
			{8'd55, 8'd127}: color_data = 12'he00;
			{8'd55, 8'd128}: color_data = 12'he00;
			{8'd55, 8'd129}: color_data = 12'he00;
			{8'd55, 8'd130}: color_data = 12'he00;
			{8'd55, 8'd131}: color_data = 12'he00;
			{8'd55, 8'd132}: color_data = 12'he00;
			{8'd55, 8'd133}: color_data = 12'he00;
			{8'd55, 8'd138}: color_data = 12'he00;
			{8'd55, 8'd139}: color_data = 12'he00;
			{8'd55, 8'd140}: color_data = 12'he00;
			{8'd55, 8'd141}: color_data = 12'he00;
			{8'd55, 8'd142}: color_data = 12'he00;
			{8'd55, 8'd143}: color_data = 12'he01;
			{8'd55, 8'd144}: color_data = 12'he00;
			{8'd56, 8'd3}: color_data = 12'h000;
			{8'd56, 8'd4}: color_data = 12'h000;
			{8'd56, 8'd5}: color_data = 12'h540;
			{8'd56, 8'd6}: color_data = 12'hfd0;
			{8'd56, 8'd7}: color_data = 12'hfd0;
			{8'd56, 8'd8}: color_data = 12'hfd0;
			{8'd56, 8'd9}: color_data = 12'hfd0;
			{8'd56, 8'd10}: color_data = 12'hfc0;
			{8'd56, 8'd11}: color_data = 12'hfc0;
			{8'd56, 8'd12}: color_data = 12'hfc0;
			{8'd56, 8'd13}: color_data = 12'hfc0;
			{8'd56, 8'd14}: color_data = 12'hfc0;
			{8'd56, 8'd15}: color_data = 12'hfc0;
			{8'd56, 8'd16}: color_data = 12'hfc0;
			{8'd56, 8'd17}: color_data = 12'hfc0;
			{8'd56, 8'd18}: color_data = 12'hfc0;
			{8'd56, 8'd19}: color_data = 12'hfc0;
			{8'd56, 8'd20}: color_data = 12'hfc0;
			{8'd56, 8'd21}: color_data = 12'hfc0;
			{8'd56, 8'd22}: color_data = 12'hfc0;
			{8'd56, 8'd23}: color_data = 12'hfc0;
			{8'd56, 8'd24}: color_data = 12'hfc0;
			{8'd56, 8'd25}: color_data = 12'hfc0;
			{8'd56, 8'd26}: color_data = 12'hfd0;
			{8'd56, 8'd27}: color_data = 12'hdb0;
			{8'd56, 8'd28}: color_data = 12'h220;
			{8'd56, 8'd29}: color_data = 12'h000;
			{8'd56, 8'd30}: color_data = 12'h000;
			{8'd56, 8'd31}: color_data = 12'h000;
			{8'd56, 8'd32}: color_data = 12'h000;
			{8'd56, 8'd33}: color_data = 12'h000;
			{8'd56, 8'd34}: color_data = 12'h000;
			{8'd56, 8'd35}: color_data = 12'h020;
			{8'd56, 8'd36}: color_data = 12'h141;
			{8'd56, 8'd37}: color_data = 12'h372;
			{8'd56, 8'd38}: color_data = 12'h3a3;
			{8'd56, 8'd39}: color_data = 12'h4b3;
			{8'd56, 8'd40}: color_data = 12'h4b3;
			{8'd56, 8'd41}: color_data = 12'h4b3;
			{8'd56, 8'd42}: color_data = 12'h4b3;
			{8'd56, 8'd43}: color_data = 12'h4a3;
			{8'd56, 8'd44}: color_data = 12'h4a3;
			{8'd56, 8'd45}: color_data = 12'h4a3;
			{8'd56, 8'd46}: color_data = 12'h4a3;
			{8'd56, 8'd47}: color_data = 12'h4a3;
			{8'd56, 8'd48}: color_data = 12'h4a3;
			{8'd56, 8'd49}: color_data = 12'h4a3;
			{8'd56, 8'd50}: color_data = 12'h4a3;
			{8'd56, 8'd51}: color_data = 12'h4a3;
			{8'd56, 8'd52}: color_data = 12'h4a3;
			{8'd56, 8'd53}: color_data = 12'h4a3;
			{8'd56, 8'd54}: color_data = 12'h4a3;
			{8'd56, 8'd55}: color_data = 12'h4a3;
			{8'd56, 8'd56}: color_data = 12'h4a3;
			{8'd56, 8'd57}: color_data = 12'h4a3;
			{8'd56, 8'd58}: color_data = 12'h4a3;
			{8'd56, 8'd59}: color_data = 12'h4a3;
			{8'd56, 8'd60}: color_data = 12'h4a3;
			{8'd56, 8'd61}: color_data = 12'h4a3;
			{8'd56, 8'd62}: color_data = 12'h4b3;
			{8'd56, 8'd63}: color_data = 12'h4b3;
			{8'd56, 8'd64}: color_data = 12'h4b3;
			{8'd56, 8'd65}: color_data = 12'h4b3;
			{8'd56, 8'd66}: color_data = 12'h4b3;
			{8'd56, 8'd67}: color_data = 12'h382;
			{8'd56, 8'd68}: color_data = 12'h000;
			{8'd56, 8'd69}: color_data = 12'h000;
			{8'd56, 8'd70}: color_data = 12'h000;
			{8'd56, 8'd71}: color_data = 12'h000;
			{8'd56, 8'd72}: color_data = 12'h000;
			{8'd56, 8'd73}: color_data = 12'h000;
			{8'd56, 8'd74}: color_data = 12'h000;
			{8'd56, 8'd100}: color_data = 12'he00;
			{8'd56, 8'd101}: color_data = 12'hf01;
			{8'd56, 8'd102}: color_data = 12'he00;
			{8'd56, 8'd103}: color_data = 12'he00;
			{8'd56, 8'd104}: color_data = 12'he00;
			{8'd56, 8'd105}: color_data = 12'he00;
			{8'd56, 8'd106}: color_data = 12'hc00;
			{8'd56, 8'd111}: color_data = 12'he00;
			{8'd56, 8'd112}: color_data = 12'he01;
			{8'd56, 8'd113}: color_data = 12'hf01;
			{8'd56, 8'd114}: color_data = 12'hf01;
			{8'd56, 8'd115}: color_data = 12'he01;
			{8'd56, 8'd116}: color_data = 12'he01;
			{8'd56, 8'd117}: color_data = 12'he01;
			{8'd56, 8'd118}: color_data = 12'he01;
			{8'd56, 8'd119}: color_data = 12'hf01;
			{8'd56, 8'd120}: color_data = 12'hf01;
			{8'd56, 8'd121}: color_data = 12'hf01;
			{8'd56, 8'd122}: color_data = 12'hf01;
			{8'd56, 8'd123}: color_data = 12'hf01;
			{8'd56, 8'd124}: color_data = 12'hf01;
			{8'd56, 8'd125}: color_data = 12'hf01;
			{8'd56, 8'd126}: color_data = 12'hf01;
			{8'd56, 8'd127}: color_data = 12'hf01;
			{8'd56, 8'd128}: color_data = 12'hf01;
			{8'd56, 8'd129}: color_data = 12'hf01;
			{8'd56, 8'd130}: color_data = 12'hf01;
			{8'd56, 8'd131}: color_data = 12'hf01;
			{8'd56, 8'd132}: color_data = 12'hf01;
			{8'd56, 8'd133}: color_data = 12'he00;
			{8'd56, 8'd138}: color_data = 12'he00;
			{8'd56, 8'd139}: color_data = 12'he00;
			{8'd56, 8'd140}: color_data = 12'he00;
			{8'd56, 8'd141}: color_data = 12'he00;
			{8'd56, 8'd142}: color_data = 12'he00;
			{8'd56, 8'd143}: color_data = 12'he01;
			{8'd56, 8'd144}: color_data = 12'he00;
			{8'd57, 8'd3}: color_data = 12'h000;
			{8'd57, 8'd4}: color_data = 12'h000;
			{8'd57, 8'd5}: color_data = 12'h330;
			{8'd57, 8'd6}: color_data = 12'hfd0;
			{8'd57, 8'd7}: color_data = 12'hfd0;
			{8'd57, 8'd8}: color_data = 12'hfc0;
			{8'd57, 8'd9}: color_data = 12'hfc0;
			{8'd57, 8'd10}: color_data = 12'hfc0;
			{8'd57, 8'd11}: color_data = 12'hfc0;
			{8'd57, 8'd12}: color_data = 12'hfc0;
			{8'd57, 8'd13}: color_data = 12'hfc0;
			{8'd57, 8'd14}: color_data = 12'hfc0;
			{8'd57, 8'd15}: color_data = 12'hfc0;
			{8'd57, 8'd16}: color_data = 12'hfc0;
			{8'd57, 8'd17}: color_data = 12'hfc0;
			{8'd57, 8'd18}: color_data = 12'hfc0;
			{8'd57, 8'd19}: color_data = 12'hfc0;
			{8'd57, 8'd20}: color_data = 12'hfc0;
			{8'd57, 8'd21}: color_data = 12'hfc0;
			{8'd57, 8'd22}: color_data = 12'hfc0;
			{8'd57, 8'd23}: color_data = 12'hfc0;
			{8'd57, 8'd24}: color_data = 12'hfc0;
			{8'd57, 8'd25}: color_data = 12'hfc0;
			{8'd57, 8'd26}: color_data = 12'hfc0;
			{8'd57, 8'd27}: color_data = 12'hfd0;
			{8'd57, 8'd28}: color_data = 12'hca0;
			{8'd57, 8'd29}: color_data = 12'h110;
			{8'd57, 8'd30}: color_data = 12'h000;
			{8'd57, 8'd31}: color_data = 12'h000;
			{8'd57, 8'd32}: color_data = 12'h000;
			{8'd57, 8'd33}: color_data = 12'h000;
			{8'd57, 8'd34}: color_data = 12'h131;
			{8'd57, 8'd35}: color_data = 12'h4b3;
			{8'd57, 8'd36}: color_data = 12'h4b3;
			{8'd57, 8'd37}: color_data = 12'h4b3;
			{8'd57, 8'd38}: color_data = 12'h4b3;
			{8'd57, 8'd39}: color_data = 12'h4a3;
			{8'd57, 8'd40}: color_data = 12'h4a3;
			{8'd57, 8'd41}: color_data = 12'h4a3;
			{8'd57, 8'd42}: color_data = 12'h4a3;
			{8'd57, 8'd43}: color_data = 12'h4a3;
			{8'd57, 8'd44}: color_data = 12'h4a3;
			{8'd57, 8'd45}: color_data = 12'h4a3;
			{8'd57, 8'd46}: color_data = 12'h4a3;
			{8'd57, 8'd47}: color_data = 12'h4a3;
			{8'd57, 8'd48}: color_data = 12'h4a3;
			{8'd57, 8'd49}: color_data = 12'h4a3;
			{8'd57, 8'd50}: color_data = 12'h4a3;
			{8'd57, 8'd51}: color_data = 12'h4a3;
			{8'd57, 8'd52}: color_data = 12'h4a3;
			{8'd57, 8'd53}: color_data = 12'h4a3;
			{8'd57, 8'd54}: color_data = 12'h4a3;
			{8'd57, 8'd55}: color_data = 12'h4a3;
			{8'd57, 8'd56}: color_data = 12'h4a3;
			{8'd57, 8'd57}: color_data = 12'h4a3;
			{8'd57, 8'd58}: color_data = 12'h4a3;
			{8'd57, 8'd59}: color_data = 12'h4a3;
			{8'd57, 8'd60}: color_data = 12'h4a3;
			{8'd57, 8'd61}: color_data = 12'h4a3;
			{8'd57, 8'd62}: color_data = 12'h4a3;
			{8'd57, 8'd63}: color_data = 12'h4a3;
			{8'd57, 8'd64}: color_data = 12'h4a3;
			{8'd57, 8'd65}: color_data = 12'h4a3;
			{8'd57, 8'd66}: color_data = 12'h4b3;
			{8'd57, 8'd67}: color_data = 12'h3a3;
			{8'd57, 8'd68}: color_data = 12'h000;
			{8'd57, 8'd69}: color_data = 12'h000;
			{8'd57, 8'd70}: color_data = 12'h000;
			{8'd57, 8'd71}: color_data = 12'h000;
			{8'd57, 8'd72}: color_data = 12'h000;
			{8'd57, 8'd73}: color_data = 12'h000;
			{8'd57, 8'd74}: color_data = 12'h000;
			{8'd57, 8'd100}: color_data = 12'he00;
			{8'd57, 8'd101}: color_data = 12'hf01;
			{8'd57, 8'd102}: color_data = 12'he00;
			{8'd57, 8'd103}: color_data = 12'he00;
			{8'd57, 8'd104}: color_data = 12'he00;
			{8'd57, 8'd105}: color_data = 12'he00;
			{8'd57, 8'd106}: color_data = 12'hc00;
			{8'd57, 8'd111}: color_data = 12'he01;
			{8'd57, 8'd112}: color_data = 12'he00;
			{8'd57, 8'd113}: color_data = 12'he00;
			{8'd57, 8'd114}: color_data = 12'he00;
			{8'd57, 8'd115}: color_data = 12'he00;
			{8'd57, 8'd116}: color_data = 12'he01;
			{8'd57, 8'd117}: color_data = 12'he01;
			{8'd57, 8'd118}: color_data = 12'he00;
			{8'd57, 8'd119}: color_data = 12'he00;
			{8'd57, 8'd120}: color_data = 12'he00;
			{8'd57, 8'd121}: color_data = 12'he00;
			{8'd57, 8'd122}: color_data = 12'he00;
			{8'd57, 8'd123}: color_data = 12'he00;
			{8'd57, 8'd124}: color_data = 12'he00;
			{8'd57, 8'd125}: color_data = 12'he00;
			{8'd57, 8'd126}: color_data = 12'he00;
			{8'd57, 8'd127}: color_data = 12'he00;
			{8'd57, 8'd128}: color_data = 12'he00;
			{8'd57, 8'd129}: color_data = 12'he00;
			{8'd57, 8'd130}: color_data = 12'he00;
			{8'd57, 8'd131}: color_data = 12'he00;
			{8'd57, 8'd132}: color_data = 12'hf01;
			{8'd57, 8'd133}: color_data = 12'he00;
			{8'd57, 8'd138}: color_data = 12'he00;
			{8'd57, 8'd139}: color_data = 12'he00;
			{8'd57, 8'd140}: color_data = 12'he00;
			{8'd57, 8'd141}: color_data = 12'he00;
			{8'd57, 8'd142}: color_data = 12'he00;
			{8'd57, 8'd143}: color_data = 12'he01;
			{8'd57, 8'd144}: color_data = 12'he00;
			{8'd58, 8'd3}: color_data = 12'h000;
			{8'd58, 8'd4}: color_data = 12'h000;
			{8'd58, 8'd5}: color_data = 12'h220;
			{8'd58, 8'd6}: color_data = 12'hfc0;
			{8'd58, 8'd7}: color_data = 12'hfd0;
			{8'd58, 8'd8}: color_data = 12'hfc0;
			{8'd58, 8'd9}: color_data = 12'hfc0;
			{8'd58, 8'd10}: color_data = 12'hfc0;
			{8'd58, 8'd11}: color_data = 12'hfc0;
			{8'd58, 8'd12}: color_data = 12'hfc0;
			{8'd58, 8'd13}: color_data = 12'hfc0;
			{8'd58, 8'd14}: color_data = 12'hfc0;
			{8'd58, 8'd15}: color_data = 12'hfc0;
			{8'd58, 8'd16}: color_data = 12'hfc0;
			{8'd58, 8'd17}: color_data = 12'hfc0;
			{8'd58, 8'd18}: color_data = 12'hfc0;
			{8'd58, 8'd19}: color_data = 12'hfc0;
			{8'd58, 8'd20}: color_data = 12'hfc0;
			{8'd58, 8'd21}: color_data = 12'hfc0;
			{8'd58, 8'd22}: color_data = 12'hfc0;
			{8'd58, 8'd23}: color_data = 12'hfc0;
			{8'd58, 8'd24}: color_data = 12'hfc0;
			{8'd58, 8'd25}: color_data = 12'hfc0;
			{8'd58, 8'd26}: color_data = 12'hfc0;
			{8'd58, 8'd27}: color_data = 12'hfc0;
			{8'd58, 8'd28}: color_data = 12'hfd0;
			{8'd58, 8'd29}: color_data = 12'hb90;
			{8'd58, 8'd30}: color_data = 12'h000;
			{8'd58, 8'd31}: color_data = 12'h000;
			{8'd58, 8'd32}: color_data = 12'h000;
			{8'd58, 8'd33}: color_data = 12'h000;
			{8'd58, 8'd34}: color_data = 12'h141;
			{8'd58, 8'd35}: color_data = 12'h4b3;
			{8'd58, 8'd36}: color_data = 12'h4a3;
			{8'd58, 8'd37}: color_data = 12'h4a3;
			{8'd58, 8'd38}: color_data = 12'h4a3;
			{8'd58, 8'd39}: color_data = 12'h4a3;
			{8'd58, 8'd40}: color_data = 12'h4a3;
			{8'd58, 8'd41}: color_data = 12'h4a3;
			{8'd58, 8'd42}: color_data = 12'h4a3;
			{8'd58, 8'd43}: color_data = 12'h4a3;
			{8'd58, 8'd44}: color_data = 12'h4a3;
			{8'd58, 8'd45}: color_data = 12'h4a3;
			{8'd58, 8'd46}: color_data = 12'h4a3;
			{8'd58, 8'd47}: color_data = 12'h4a3;
			{8'd58, 8'd48}: color_data = 12'h4a3;
			{8'd58, 8'd49}: color_data = 12'h4a3;
			{8'd58, 8'd50}: color_data = 12'h4a3;
			{8'd58, 8'd51}: color_data = 12'h4a3;
			{8'd58, 8'd52}: color_data = 12'h4a3;
			{8'd58, 8'd53}: color_data = 12'h4a3;
			{8'd58, 8'd54}: color_data = 12'h4a3;
			{8'd58, 8'd55}: color_data = 12'h4a3;
			{8'd58, 8'd56}: color_data = 12'h4a3;
			{8'd58, 8'd57}: color_data = 12'h4a3;
			{8'd58, 8'd58}: color_data = 12'h4a3;
			{8'd58, 8'd59}: color_data = 12'h4a3;
			{8'd58, 8'd60}: color_data = 12'h4a3;
			{8'd58, 8'd61}: color_data = 12'h4a3;
			{8'd58, 8'd62}: color_data = 12'h4a3;
			{8'd58, 8'd63}: color_data = 12'h4b3;
			{8'd58, 8'd64}: color_data = 12'h4b3;
			{8'd58, 8'd65}: color_data = 12'h4b3;
			{8'd58, 8'd66}: color_data = 12'h4b3;
			{8'd58, 8'd67}: color_data = 12'h4b3;
			{8'd58, 8'd68}: color_data = 12'h020;
			{8'd58, 8'd69}: color_data = 12'h000;
			{8'd58, 8'd70}: color_data = 12'h000;
			{8'd58, 8'd71}: color_data = 12'h000;
			{8'd58, 8'd72}: color_data = 12'h000;
			{8'd58, 8'd73}: color_data = 12'h000;
			{8'd58, 8'd74}: color_data = 12'h000;
			{8'd58, 8'd75}: color_data = 12'h000;
			{8'd58, 8'd100}: color_data = 12'he00;
			{8'd58, 8'd101}: color_data = 12'hf01;
			{8'd58, 8'd102}: color_data = 12'he00;
			{8'd58, 8'd103}: color_data = 12'he00;
			{8'd58, 8'd104}: color_data = 12'he00;
			{8'd58, 8'd105}: color_data = 12'he00;
			{8'd58, 8'd106}: color_data = 12'hc00;
			{8'd58, 8'd111}: color_data = 12'he01;
			{8'd58, 8'd112}: color_data = 12'he00;
			{8'd58, 8'd113}: color_data = 12'he00;
			{8'd58, 8'd114}: color_data = 12'he00;
			{8'd58, 8'd115}: color_data = 12'he00;
			{8'd58, 8'd116}: color_data = 12'he01;
			{8'd58, 8'd117}: color_data = 12'he01;
			{8'd58, 8'd118}: color_data = 12'he00;
			{8'd58, 8'd119}: color_data = 12'he00;
			{8'd58, 8'd120}: color_data = 12'he00;
			{8'd58, 8'd121}: color_data = 12'he00;
			{8'd58, 8'd122}: color_data = 12'he00;
			{8'd58, 8'd123}: color_data = 12'he00;
			{8'd58, 8'd124}: color_data = 12'he00;
			{8'd58, 8'd125}: color_data = 12'he00;
			{8'd58, 8'd126}: color_data = 12'he00;
			{8'd58, 8'd127}: color_data = 12'he00;
			{8'd58, 8'd128}: color_data = 12'he00;
			{8'd58, 8'd129}: color_data = 12'he00;
			{8'd58, 8'd130}: color_data = 12'he00;
			{8'd58, 8'd131}: color_data = 12'he00;
			{8'd58, 8'd132}: color_data = 12'hf01;
			{8'd58, 8'd133}: color_data = 12'he00;
			{8'd58, 8'd138}: color_data = 12'he00;
			{8'd58, 8'd139}: color_data = 12'he00;
			{8'd58, 8'd140}: color_data = 12'he00;
			{8'd58, 8'd141}: color_data = 12'he00;
			{8'd58, 8'd142}: color_data = 12'he00;
			{8'd58, 8'd143}: color_data = 12'he01;
			{8'd58, 8'd144}: color_data = 12'he00;
			{8'd59, 8'd3}: color_data = 12'h000;
			{8'd59, 8'd4}: color_data = 12'h000;
			{8'd59, 8'd5}: color_data = 12'h110;
			{8'd59, 8'd6}: color_data = 12'hec0;
			{8'd59, 8'd7}: color_data = 12'hfd0;
			{8'd59, 8'd8}: color_data = 12'hfc0;
			{8'd59, 8'd9}: color_data = 12'hfc0;
			{8'd59, 8'd10}: color_data = 12'hfc0;
			{8'd59, 8'd11}: color_data = 12'hfc0;
			{8'd59, 8'd12}: color_data = 12'hfc0;
			{8'd59, 8'd13}: color_data = 12'hfc0;
			{8'd59, 8'd14}: color_data = 12'hfc0;
			{8'd59, 8'd15}: color_data = 12'hfc0;
			{8'd59, 8'd16}: color_data = 12'hfc0;
			{8'd59, 8'd17}: color_data = 12'hfc0;
			{8'd59, 8'd18}: color_data = 12'hfc0;
			{8'd59, 8'd19}: color_data = 12'hfc0;
			{8'd59, 8'd20}: color_data = 12'hfc0;
			{8'd59, 8'd21}: color_data = 12'hfc0;
			{8'd59, 8'd22}: color_data = 12'hfc0;
			{8'd59, 8'd23}: color_data = 12'hfc0;
			{8'd59, 8'd24}: color_data = 12'hfc0;
			{8'd59, 8'd25}: color_data = 12'hfc0;
			{8'd59, 8'd26}: color_data = 12'hfc0;
			{8'd59, 8'd27}: color_data = 12'hfc0;
			{8'd59, 8'd28}: color_data = 12'hfd0;
			{8'd59, 8'd29}: color_data = 12'heb0;
			{8'd59, 8'd30}: color_data = 12'h100;
			{8'd59, 8'd31}: color_data = 12'h000;
			{8'd59, 8'd32}: color_data = 12'h000;
			{8'd59, 8'd33}: color_data = 12'h000;
			{8'd59, 8'd34}: color_data = 12'h120;
			{8'd59, 8'd35}: color_data = 12'h4b3;
			{8'd59, 8'd36}: color_data = 12'h4a3;
			{8'd59, 8'd37}: color_data = 12'h4a3;
			{8'd59, 8'd38}: color_data = 12'h4a3;
			{8'd59, 8'd39}: color_data = 12'h4a3;
			{8'd59, 8'd40}: color_data = 12'h4a3;
			{8'd59, 8'd41}: color_data = 12'h4a3;
			{8'd59, 8'd42}: color_data = 12'h4a3;
			{8'd59, 8'd43}: color_data = 12'h4a3;
			{8'd59, 8'd44}: color_data = 12'h4a3;
			{8'd59, 8'd45}: color_data = 12'h4a3;
			{8'd59, 8'd46}: color_data = 12'h4a3;
			{8'd59, 8'd47}: color_data = 12'h4a3;
			{8'd59, 8'd48}: color_data = 12'h4a3;
			{8'd59, 8'd49}: color_data = 12'h4a3;
			{8'd59, 8'd50}: color_data = 12'h4a3;
			{8'd59, 8'd51}: color_data = 12'h4a3;
			{8'd59, 8'd52}: color_data = 12'h4a3;
			{8'd59, 8'd53}: color_data = 12'h4a3;
			{8'd59, 8'd54}: color_data = 12'h4a3;
			{8'd59, 8'd55}: color_data = 12'h4a3;
			{8'd59, 8'd56}: color_data = 12'h4a3;
			{8'd59, 8'd57}: color_data = 12'h4a3;
			{8'd59, 8'd58}: color_data = 12'h4a3;
			{8'd59, 8'd59}: color_data = 12'h4a3;
			{8'd59, 8'd60}: color_data = 12'h4a3;
			{8'd59, 8'd61}: color_data = 12'h4b3;
			{8'd59, 8'd62}: color_data = 12'h4b3;
			{8'd59, 8'd63}: color_data = 12'h4a3;
			{8'd59, 8'd64}: color_data = 12'h392;
			{8'd59, 8'd65}: color_data = 12'h372;
			{8'd59, 8'd66}: color_data = 12'h261;
			{8'd59, 8'd67}: color_data = 12'h141;
			{8'd59, 8'd68}: color_data = 12'h000;
			{8'd59, 8'd69}: color_data = 12'h000;
			{8'd59, 8'd70}: color_data = 12'h000;
			{8'd59, 8'd71}: color_data = 12'h000;
			{8'd59, 8'd72}: color_data = 12'h000;
			{8'd59, 8'd73}: color_data = 12'h000;
			{8'd59, 8'd74}: color_data = 12'h000;
			{8'd59, 8'd75}: color_data = 12'h000;
			{8'd59, 8'd100}: color_data = 12'he00;
			{8'd59, 8'd101}: color_data = 12'hf01;
			{8'd59, 8'd102}: color_data = 12'he00;
			{8'd59, 8'd103}: color_data = 12'he00;
			{8'd59, 8'd104}: color_data = 12'he00;
			{8'd59, 8'd105}: color_data = 12'he00;
			{8'd59, 8'd106}: color_data = 12'hc00;
			{8'd59, 8'd111}: color_data = 12'he01;
			{8'd59, 8'd112}: color_data = 12'he00;
			{8'd59, 8'd113}: color_data = 12'he00;
			{8'd59, 8'd114}: color_data = 12'he00;
			{8'd59, 8'd115}: color_data = 12'he00;
			{8'd59, 8'd116}: color_data = 12'he01;
			{8'd59, 8'd117}: color_data = 12'he01;
			{8'd59, 8'd118}: color_data = 12'he00;
			{8'd59, 8'd119}: color_data = 12'he00;
			{8'd59, 8'd120}: color_data = 12'he00;
			{8'd59, 8'd121}: color_data = 12'he00;
			{8'd59, 8'd122}: color_data = 12'he00;
			{8'd59, 8'd123}: color_data = 12'he00;
			{8'd59, 8'd124}: color_data = 12'he00;
			{8'd59, 8'd125}: color_data = 12'he00;
			{8'd59, 8'd126}: color_data = 12'he00;
			{8'd59, 8'd127}: color_data = 12'he00;
			{8'd59, 8'd128}: color_data = 12'he00;
			{8'd59, 8'd129}: color_data = 12'he00;
			{8'd59, 8'd130}: color_data = 12'he00;
			{8'd59, 8'd131}: color_data = 12'he00;
			{8'd59, 8'd132}: color_data = 12'hf01;
			{8'd59, 8'd133}: color_data = 12'he00;
			{8'd59, 8'd138}: color_data = 12'he00;
			{8'd59, 8'd139}: color_data = 12'he00;
			{8'd59, 8'd140}: color_data = 12'he00;
			{8'd59, 8'd141}: color_data = 12'he00;
			{8'd59, 8'd142}: color_data = 12'he00;
			{8'd59, 8'd143}: color_data = 12'he01;
			{8'd59, 8'd144}: color_data = 12'he00;
			{8'd60, 8'd3}: color_data = 12'h000;
			{8'd60, 8'd4}: color_data = 12'h000;
			{8'd60, 8'd5}: color_data = 12'h000;
			{8'd60, 8'd6}: color_data = 12'hdb0;
			{8'd60, 8'd7}: color_data = 12'hfd0;
			{8'd60, 8'd8}: color_data = 12'hfc0;
			{8'd60, 8'd9}: color_data = 12'hfc0;
			{8'd60, 8'd10}: color_data = 12'hfc0;
			{8'd60, 8'd11}: color_data = 12'hfc0;
			{8'd60, 8'd12}: color_data = 12'hfc0;
			{8'd60, 8'd13}: color_data = 12'hfc0;
			{8'd60, 8'd14}: color_data = 12'hfc0;
			{8'd60, 8'd15}: color_data = 12'hfc0;
			{8'd60, 8'd16}: color_data = 12'hfc0;
			{8'd60, 8'd17}: color_data = 12'hfd0;
			{8'd60, 8'd18}: color_data = 12'hfd0;
			{8'd60, 8'd19}: color_data = 12'hfd0;
			{8'd60, 8'd20}: color_data = 12'hfd0;
			{8'd60, 8'd21}: color_data = 12'hfd0;
			{8'd60, 8'd22}: color_data = 12'hfd0;
			{8'd60, 8'd23}: color_data = 12'hfc0;
			{8'd60, 8'd24}: color_data = 12'hfc0;
			{8'd60, 8'd25}: color_data = 12'hfc0;
			{8'd60, 8'd26}: color_data = 12'hfc0;
			{8'd60, 8'd27}: color_data = 12'hfc0;
			{8'd60, 8'd28}: color_data = 12'hfd0;
			{8'd60, 8'd29}: color_data = 12'heb0;
			{8'd60, 8'd30}: color_data = 12'h110;
			{8'd60, 8'd31}: color_data = 12'h000;
			{8'd60, 8'd32}: color_data = 12'h000;
			{8'd60, 8'd33}: color_data = 12'h000;
			{8'd60, 8'd34}: color_data = 12'h020;
			{8'd60, 8'd35}: color_data = 12'h4a3;
			{8'd60, 8'd36}: color_data = 12'h4b3;
			{8'd60, 8'd37}: color_data = 12'h4a3;
			{8'd60, 8'd38}: color_data = 12'h4a3;
			{8'd60, 8'd39}: color_data = 12'h4a3;
			{8'd60, 8'd40}: color_data = 12'h4a3;
			{8'd60, 8'd41}: color_data = 12'h4a3;
			{8'd60, 8'd42}: color_data = 12'h4a3;
			{8'd60, 8'd43}: color_data = 12'h4a3;
			{8'd60, 8'd44}: color_data = 12'h4a3;
			{8'd60, 8'd45}: color_data = 12'h4a3;
			{8'd60, 8'd46}: color_data = 12'h4a3;
			{8'd60, 8'd47}: color_data = 12'h4a3;
			{8'd60, 8'd48}: color_data = 12'h4a3;
			{8'd60, 8'd49}: color_data = 12'h4a3;
			{8'd60, 8'd50}: color_data = 12'h4a3;
			{8'd60, 8'd51}: color_data = 12'h4b3;
			{8'd60, 8'd52}: color_data = 12'h4b3;
			{8'd60, 8'd53}: color_data = 12'h4b3;
			{8'd60, 8'd54}: color_data = 12'h4a3;
			{8'd60, 8'd55}: color_data = 12'h4a3;
			{8'd60, 8'd56}: color_data = 12'h4a3;
			{8'd60, 8'd57}: color_data = 12'h4a3;
			{8'd60, 8'd58}: color_data = 12'h4a3;
			{8'd60, 8'd59}: color_data = 12'h4a3;
			{8'd60, 8'd60}: color_data = 12'h4b3;
			{8'd60, 8'd61}: color_data = 12'h272;
			{8'd60, 8'd62}: color_data = 12'h120;
			{8'd60, 8'd63}: color_data = 12'h010;
			{8'd60, 8'd64}: color_data = 12'h000;
			{8'd60, 8'd65}: color_data = 12'h000;
			{8'd60, 8'd66}: color_data = 12'h000;
			{8'd60, 8'd67}: color_data = 12'h000;
			{8'd60, 8'd68}: color_data = 12'h000;
			{8'd60, 8'd69}: color_data = 12'h000;
			{8'd60, 8'd70}: color_data = 12'h000;
			{8'd60, 8'd71}: color_data = 12'h000;
			{8'd60, 8'd72}: color_data = 12'h000;
			{8'd60, 8'd73}: color_data = 12'h000;
			{8'd60, 8'd74}: color_data = 12'h000;
			{8'd60, 8'd75}: color_data = 12'h000;
			{8'd60, 8'd100}: color_data = 12'he00;
			{8'd60, 8'd101}: color_data = 12'hf01;
			{8'd60, 8'd102}: color_data = 12'he00;
			{8'd60, 8'd103}: color_data = 12'he00;
			{8'd60, 8'd104}: color_data = 12'he00;
			{8'd60, 8'd105}: color_data = 12'he00;
			{8'd60, 8'd106}: color_data = 12'hc00;
			{8'd60, 8'd111}: color_data = 12'he00;
			{8'd60, 8'd112}: color_data = 12'he01;
			{8'd60, 8'd113}: color_data = 12'hf01;
			{8'd60, 8'd114}: color_data = 12'hf01;
			{8'd60, 8'd115}: color_data = 12'he00;
			{8'd60, 8'd116}: color_data = 12'hd01;
			{8'd60, 8'd117}: color_data = 12'he01;
			{8'd60, 8'd118}: color_data = 12'he01;
			{8'd60, 8'd119}: color_data = 12'hf01;
			{8'd60, 8'd120}: color_data = 12'he01;
			{8'd60, 8'd121}: color_data = 12'he01;
			{8'd60, 8'd122}: color_data = 12'he01;
			{8'd60, 8'd123}: color_data = 12'he01;
			{8'd60, 8'd124}: color_data = 12'he01;
			{8'd60, 8'd125}: color_data = 12'he01;
			{8'd60, 8'd126}: color_data = 12'he01;
			{8'd60, 8'd127}: color_data = 12'he01;
			{8'd60, 8'd128}: color_data = 12'he01;
			{8'd60, 8'd129}: color_data = 12'he01;
			{8'd60, 8'd130}: color_data = 12'he01;
			{8'd60, 8'd131}: color_data = 12'he01;
			{8'd60, 8'd132}: color_data = 12'hf01;
			{8'd60, 8'd133}: color_data = 12'he00;
			{8'd60, 8'd138}: color_data = 12'he00;
			{8'd60, 8'd139}: color_data = 12'he00;
			{8'd60, 8'd140}: color_data = 12'he00;
			{8'd60, 8'd141}: color_data = 12'he00;
			{8'd60, 8'd142}: color_data = 12'he00;
			{8'd60, 8'd143}: color_data = 12'he01;
			{8'd60, 8'd144}: color_data = 12'he00;
			{8'd61, 8'd3}: color_data = 12'h000;
			{8'd61, 8'd4}: color_data = 12'h000;
			{8'd61, 8'd5}: color_data = 12'h000;
			{8'd61, 8'd6}: color_data = 12'hca0;
			{8'd61, 8'd7}: color_data = 12'hfd0;
			{8'd61, 8'd8}: color_data = 12'hfc0;
			{8'd61, 8'd9}: color_data = 12'hfc0;
			{8'd61, 8'd10}: color_data = 12'hfc0;
			{8'd61, 8'd11}: color_data = 12'hfd0;
			{8'd61, 8'd12}: color_data = 12'hfd0;
			{8'd61, 8'd13}: color_data = 12'hfd0;
			{8'd61, 8'd14}: color_data = 12'hfd0;
			{8'd61, 8'd15}: color_data = 12'hfd0;
			{8'd61, 8'd16}: color_data = 12'hfd0;
			{8'd61, 8'd17}: color_data = 12'hfc0;
			{8'd61, 8'd18}: color_data = 12'heb0;
			{8'd61, 8'd19}: color_data = 12'hca0;
			{8'd61, 8'd20}: color_data = 12'ha80;
			{8'd61, 8'd21}: color_data = 12'h760;
			{8'd61, 8'd22}: color_data = 12'h980;
			{8'd61, 8'd23}: color_data = 12'hfd0;
			{8'd61, 8'd24}: color_data = 12'hfc0;
			{8'd61, 8'd25}: color_data = 12'hfc0;
			{8'd61, 8'd26}: color_data = 12'hfc0;
			{8'd61, 8'd27}: color_data = 12'hfc0;
			{8'd61, 8'd28}: color_data = 12'hfd0;
			{8'd61, 8'd29}: color_data = 12'hec0;
			{8'd61, 8'd30}: color_data = 12'h110;
			{8'd61, 8'd31}: color_data = 12'h000;
			{8'd61, 8'd32}: color_data = 12'h000;
			{8'd61, 8'd33}: color_data = 12'h000;
			{8'd61, 8'd34}: color_data = 12'h010;
			{8'd61, 8'd35}: color_data = 12'h4a3;
			{8'd61, 8'd36}: color_data = 12'h4b3;
			{8'd61, 8'd37}: color_data = 12'h4a3;
			{8'd61, 8'd38}: color_data = 12'h4a3;
			{8'd61, 8'd39}: color_data = 12'h4a3;
			{8'd61, 8'd40}: color_data = 12'h4a3;
			{8'd61, 8'd41}: color_data = 12'h4a3;
			{8'd61, 8'd42}: color_data = 12'h4a3;
			{8'd61, 8'd43}: color_data = 12'h4a3;
			{8'd61, 8'd44}: color_data = 12'h4a3;
			{8'd61, 8'd45}: color_data = 12'h4b3;
			{8'd61, 8'd46}: color_data = 12'h4b3;
			{8'd61, 8'd47}: color_data = 12'h4b3;
			{8'd61, 8'd48}: color_data = 12'h4b3;
			{8'd61, 8'd49}: color_data = 12'h4b3;
			{8'd61, 8'd50}: color_data = 12'h4b3;
			{8'd61, 8'd51}: color_data = 12'h4a3;
			{8'd61, 8'd52}: color_data = 12'h392;
			{8'd61, 8'd53}: color_data = 12'h4a3;
			{8'd61, 8'd54}: color_data = 12'h4b3;
			{8'd61, 8'd55}: color_data = 12'h4a3;
			{8'd61, 8'd56}: color_data = 12'h4a3;
			{8'd61, 8'd57}: color_data = 12'h4a3;
			{8'd61, 8'd58}: color_data = 12'h4a3;
			{8'd61, 8'd59}: color_data = 12'h4a3;
			{8'd61, 8'd60}: color_data = 12'h4b3;
			{8'd61, 8'd61}: color_data = 12'h141;
			{8'd61, 8'd62}: color_data = 12'h000;
			{8'd61, 8'd63}: color_data = 12'h000;
			{8'd61, 8'd64}: color_data = 12'h000;
			{8'd61, 8'd65}: color_data = 12'h000;
			{8'd61, 8'd66}: color_data = 12'h000;
			{8'd61, 8'd67}: color_data = 12'h000;
			{8'd61, 8'd68}: color_data = 12'h000;
			{8'd61, 8'd69}: color_data = 12'h000;
			{8'd61, 8'd70}: color_data = 12'h000;
			{8'd61, 8'd71}: color_data = 12'h000;
			{8'd61, 8'd72}: color_data = 12'h000;
			{8'd61, 8'd73}: color_data = 12'h000;
			{8'd61, 8'd74}: color_data = 12'h000;
			{8'd61, 8'd75}: color_data = 12'h000;
			{8'd61, 8'd100}: color_data = 12'he00;
			{8'd61, 8'd101}: color_data = 12'hf01;
			{8'd61, 8'd102}: color_data = 12'he00;
			{8'd61, 8'd103}: color_data = 12'he00;
			{8'd61, 8'd104}: color_data = 12'he00;
			{8'd61, 8'd105}: color_data = 12'he00;
			{8'd61, 8'd106}: color_data = 12'hc00;
			{8'd61, 8'd111}: color_data = 12'he00;
			{8'd61, 8'd112}: color_data = 12'he00;
			{8'd61, 8'd113}: color_data = 12'he00;
			{8'd61, 8'd114}: color_data = 12'he00;
			{8'd61, 8'd115}: color_data = 12'he00;
			{8'd61, 8'd116}: color_data = 12'hd01;
			{8'd61, 8'd117}: color_data = 12'he01;
			{8'd61, 8'd118}: color_data = 12'he00;
			{8'd61, 8'd119}: color_data = 12'he00;
			{8'd61, 8'd120}: color_data = 12'he00;
			{8'd61, 8'd121}: color_data = 12'he00;
			{8'd61, 8'd122}: color_data = 12'he00;
			{8'd61, 8'd123}: color_data = 12'he00;
			{8'd61, 8'd124}: color_data = 12'he00;
			{8'd61, 8'd125}: color_data = 12'he00;
			{8'd61, 8'd126}: color_data = 12'he00;
			{8'd61, 8'd127}: color_data = 12'he00;
			{8'd61, 8'd128}: color_data = 12'he00;
			{8'd61, 8'd129}: color_data = 12'he00;
			{8'd61, 8'd130}: color_data = 12'he00;
			{8'd61, 8'd131}: color_data = 12'he00;
			{8'd61, 8'd132}: color_data = 12'he00;
			{8'd61, 8'd133}: color_data = 12'he00;
			{8'd61, 8'd138}: color_data = 12'he00;
			{8'd61, 8'd139}: color_data = 12'he00;
			{8'd61, 8'd140}: color_data = 12'he00;
			{8'd61, 8'd141}: color_data = 12'he00;
			{8'd61, 8'd142}: color_data = 12'he00;
			{8'd61, 8'd143}: color_data = 12'he01;
			{8'd61, 8'd144}: color_data = 12'he00;
			{8'd62, 8'd3}: color_data = 12'h000;
			{8'd62, 8'd4}: color_data = 12'h000;
			{8'd62, 8'd5}: color_data = 12'h000;
			{8'd62, 8'd6}: color_data = 12'hb90;
			{8'd62, 8'd7}: color_data = 12'hfd0;
			{8'd62, 8'd8}: color_data = 12'hfd0;
			{8'd62, 8'd9}: color_data = 12'hfd0;
			{8'd62, 8'd10}: color_data = 12'hfd0;
			{8'd62, 8'd11}: color_data = 12'hfc0;
			{8'd62, 8'd12}: color_data = 12'heb0;
			{8'd62, 8'd13}: color_data = 12'hca0;
			{8'd62, 8'd14}: color_data = 12'ha80;
			{8'd62, 8'd15}: color_data = 12'h760;
			{8'd62, 8'd16}: color_data = 12'h540;
			{8'd62, 8'd17}: color_data = 12'h320;
			{8'd62, 8'd18}: color_data = 12'h110;
			{8'd62, 8'd19}: color_data = 12'h000;
			{8'd62, 8'd20}: color_data = 12'h000;
			{8'd62, 8'd21}: color_data = 12'h000;
			{8'd62, 8'd22}: color_data = 12'h650;
			{8'd62, 8'd23}: color_data = 12'hfd0;
			{8'd62, 8'd24}: color_data = 12'hfc0;
			{8'd62, 8'd25}: color_data = 12'hfc0;
			{8'd62, 8'd26}: color_data = 12'hfc0;
			{8'd62, 8'd27}: color_data = 12'hfc0;
			{8'd62, 8'd28}: color_data = 12'hfd0;
			{8'd62, 8'd29}: color_data = 12'hec0;
			{8'd62, 8'd30}: color_data = 12'h110;
			{8'd62, 8'd31}: color_data = 12'h000;
			{8'd62, 8'd32}: color_data = 12'h000;
			{8'd62, 8'd33}: color_data = 12'h000;
			{8'd62, 8'd34}: color_data = 12'h000;
			{8'd62, 8'd35}: color_data = 12'h392;
			{8'd62, 8'd36}: color_data = 12'h4b3;
			{8'd62, 8'd37}: color_data = 12'h4a3;
			{8'd62, 8'd38}: color_data = 12'h4a3;
			{8'd62, 8'd39}: color_data = 12'h4a3;
			{8'd62, 8'd40}: color_data = 12'h4a3;
			{8'd62, 8'd41}: color_data = 12'h4a3;
			{8'd62, 8'd42}: color_data = 12'h4a3;
			{8'd62, 8'd43}: color_data = 12'h4a3;
			{8'd62, 8'd44}: color_data = 12'h4b3;
			{8'd62, 8'd45}: color_data = 12'h4a3;
			{8'd62, 8'd46}: color_data = 12'h392;
			{8'd62, 8'd47}: color_data = 12'h382;
			{8'd62, 8'd48}: color_data = 12'h262;
			{8'd62, 8'd49}: color_data = 12'h141;
			{8'd62, 8'd50}: color_data = 12'h130;
			{8'd62, 8'd51}: color_data = 12'h010;
			{8'd62, 8'd52}: color_data = 12'h000;
			{8'd62, 8'd53}: color_data = 12'h392;
			{8'd62, 8'd54}: color_data = 12'h4b3;
			{8'd62, 8'd55}: color_data = 12'h4a3;
			{8'd62, 8'd56}: color_data = 12'h4a3;
			{8'd62, 8'd57}: color_data = 12'h4a3;
			{8'd62, 8'd58}: color_data = 12'h4a3;
			{8'd62, 8'd59}: color_data = 12'h4b3;
			{8'd62, 8'd60}: color_data = 12'h4b3;
			{8'd62, 8'd61}: color_data = 12'h120;
			{8'd62, 8'd62}: color_data = 12'h000;
			{8'd62, 8'd63}: color_data = 12'h000;
			{8'd62, 8'd64}: color_data = 12'h000;
			{8'd62, 8'd65}: color_data = 12'h000;
			{8'd62, 8'd66}: color_data = 12'h000;
			{8'd62, 8'd67}: color_data = 12'h000;
			{8'd62, 8'd68}: color_data = 12'h000;
			{8'd62, 8'd69}: color_data = 12'h000;
			{8'd62, 8'd70}: color_data = 12'h000;
			{8'd62, 8'd71}: color_data = 12'h000;
			{8'd62, 8'd72}: color_data = 12'h000;
			{8'd62, 8'd73}: color_data = 12'h000;
			{8'd62, 8'd100}: color_data = 12'he00;
			{8'd62, 8'd101}: color_data = 12'hf01;
			{8'd62, 8'd102}: color_data = 12'he00;
			{8'd62, 8'd103}: color_data = 12'he00;
			{8'd62, 8'd104}: color_data = 12'he00;
			{8'd62, 8'd105}: color_data = 12'he00;
			{8'd62, 8'd106}: color_data = 12'hc00;
			{8'd62, 8'd138}: color_data = 12'he00;
			{8'd62, 8'd139}: color_data = 12'he00;
			{8'd62, 8'd140}: color_data = 12'he00;
			{8'd62, 8'd141}: color_data = 12'he00;
			{8'd62, 8'd142}: color_data = 12'he00;
			{8'd62, 8'd143}: color_data = 12'he01;
			{8'd62, 8'd144}: color_data = 12'he00;
			{8'd63, 8'd3}: color_data = 12'h000;
			{8'd63, 8'd4}: color_data = 12'h000;
			{8'd63, 8'd5}: color_data = 12'h000;
			{8'd63, 8'd6}: color_data = 12'h870;
			{8'd63, 8'd7}: color_data = 12'hca0;
			{8'd63, 8'd8}: color_data = 12'h980;
			{8'd63, 8'd9}: color_data = 12'h760;
			{8'd63, 8'd10}: color_data = 12'h440;
			{8'd63, 8'd11}: color_data = 12'h220;
			{8'd63, 8'd12}: color_data = 12'h100;
			{8'd63, 8'd13}: color_data = 12'h000;
			{8'd63, 8'd14}: color_data = 12'h000;
			{8'd63, 8'd15}: color_data = 12'h000;
			{8'd63, 8'd16}: color_data = 12'h000;
			{8'd63, 8'd17}: color_data = 12'h000;
			{8'd63, 8'd18}: color_data = 12'h000;
			{8'd63, 8'd19}: color_data = 12'h000;
			{8'd63, 8'd20}: color_data = 12'h000;
			{8'd63, 8'd21}: color_data = 12'h000;
			{8'd63, 8'd22}: color_data = 12'h760;
			{8'd63, 8'd23}: color_data = 12'hfd0;
			{8'd63, 8'd24}: color_data = 12'hfc0;
			{8'd63, 8'd25}: color_data = 12'hfc0;
			{8'd63, 8'd26}: color_data = 12'hfc0;
			{8'd63, 8'd27}: color_data = 12'hfc0;
			{8'd63, 8'd28}: color_data = 12'hfd0;
			{8'd63, 8'd29}: color_data = 12'hfc0;
			{8'd63, 8'd30}: color_data = 12'h210;
			{8'd63, 8'd31}: color_data = 12'h000;
			{8'd63, 8'd32}: color_data = 12'h000;
			{8'd63, 8'd33}: color_data = 12'h000;
			{8'd63, 8'd34}: color_data = 12'h000;
			{8'd63, 8'd35}: color_data = 12'h382;
			{8'd63, 8'd36}: color_data = 12'h4b3;
			{8'd63, 8'd37}: color_data = 12'h4a3;
			{8'd63, 8'd38}: color_data = 12'h4a3;
			{8'd63, 8'd39}: color_data = 12'h4a3;
			{8'd63, 8'd40}: color_data = 12'h4a3;
			{8'd63, 8'd41}: color_data = 12'h4a3;
			{8'd63, 8'd42}: color_data = 12'h4b3;
			{8'd63, 8'd43}: color_data = 12'h4a3;
			{8'd63, 8'd44}: color_data = 12'h141;
			{8'd63, 8'd45}: color_data = 12'h010;
			{8'd63, 8'd46}: color_data = 12'h000;
			{8'd63, 8'd47}: color_data = 12'h000;
			{8'd63, 8'd48}: color_data = 12'h000;
			{8'd63, 8'd49}: color_data = 12'h000;
			{8'd63, 8'd50}: color_data = 12'h000;
			{8'd63, 8'd51}: color_data = 12'h000;
			{8'd63, 8'd52}: color_data = 12'h000;
			{8'd63, 8'd53}: color_data = 12'h382;
			{8'd63, 8'd54}: color_data = 12'h4b3;
			{8'd63, 8'd55}: color_data = 12'h4a3;
			{8'd63, 8'd56}: color_data = 12'h4a3;
			{8'd63, 8'd57}: color_data = 12'h4a3;
			{8'd63, 8'd58}: color_data = 12'h4a3;
			{8'd63, 8'd59}: color_data = 12'h4b3;
			{8'd63, 8'd60}: color_data = 12'h4a3;
			{8'd63, 8'd61}: color_data = 12'h010;
			{8'd63, 8'd62}: color_data = 12'h000;
			{8'd63, 8'd63}: color_data = 12'h000;
			{8'd63, 8'd64}: color_data = 12'h000;
			{8'd63, 8'd65}: color_data = 12'h000;
			{8'd63, 8'd66}: color_data = 12'h000;
			{8'd63, 8'd67}: color_data = 12'h000;
			{8'd63, 8'd68}: color_data = 12'h000;
			{8'd63, 8'd100}: color_data = 12'he00;
			{8'd63, 8'd101}: color_data = 12'hf01;
			{8'd63, 8'd102}: color_data = 12'he00;
			{8'd63, 8'd103}: color_data = 12'he00;
			{8'd63, 8'd104}: color_data = 12'he00;
			{8'd63, 8'd105}: color_data = 12'he00;
			{8'd63, 8'd106}: color_data = 12'hc00;
			{8'd63, 8'd117}: color_data = 12'he01;
			{8'd63, 8'd118}: color_data = 12'hd00;
			{8'd63, 8'd138}: color_data = 12'he00;
			{8'd63, 8'd139}: color_data = 12'he00;
			{8'd63, 8'd140}: color_data = 12'he00;
			{8'd63, 8'd141}: color_data = 12'he00;
			{8'd63, 8'd142}: color_data = 12'he00;
			{8'd63, 8'd143}: color_data = 12'he01;
			{8'd63, 8'd144}: color_data = 12'he00;
			{8'd64, 8'd3}: color_data = 12'h000;
			{8'd64, 8'd4}: color_data = 12'h000;
			{8'd64, 8'd5}: color_data = 12'h000;
			{8'd64, 8'd6}: color_data = 12'h000;
			{8'd64, 8'd7}: color_data = 12'h000;
			{8'd64, 8'd8}: color_data = 12'h000;
			{8'd64, 8'd9}: color_data = 12'h000;
			{8'd64, 8'd10}: color_data = 12'h000;
			{8'd64, 8'd11}: color_data = 12'h000;
			{8'd64, 8'd12}: color_data = 12'h000;
			{8'd64, 8'd13}: color_data = 12'h000;
			{8'd64, 8'd14}: color_data = 12'h000;
			{8'd64, 8'd15}: color_data = 12'h000;
			{8'd64, 8'd16}: color_data = 12'h000;
			{8'd64, 8'd17}: color_data = 12'h000;
			{8'd64, 8'd18}: color_data = 12'h000;
			{8'd64, 8'd19}: color_data = 12'h000;
			{8'd64, 8'd20}: color_data = 12'h000;
			{8'd64, 8'd21}: color_data = 12'h000;
			{8'd64, 8'd22}: color_data = 12'h870;
			{8'd64, 8'd23}: color_data = 12'hfd0;
			{8'd64, 8'd24}: color_data = 12'hfc0;
			{8'd64, 8'd25}: color_data = 12'hfc0;
			{8'd64, 8'd26}: color_data = 12'hfc0;
			{8'd64, 8'd27}: color_data = 12'hfc0;
			{8'd64, 8'd28}: color_data = 12'hfd0;
			{8'd64, 8'd29}: color_data = 12'hfc0;
			{8'd64, 8'd30}: color_data = 12'h210;
			{8'd64, 8'd31}: color_data = 12'h000;
			{8'd64, 8'd32}: color_data = 12'h000;
			{8'd64, 8'd33}: color_data = 12'h000;
			{8'd64, 8'd34}: color_data = 12'h000;
			{8'd64, 8'd35}: color_data = 12'h382;
			{8'd64, 8'd36}: color_data = 12'h4b3;
			{8'd64, 8'd37}: color_data = 12'h4a3;
			{8'd64, 8'd38}: color_data = 12'h4a3;
			{8'd64, 8'd39}: color_data = 12'h4a3;
			{8'd64, 8'd40}: color_data = 12'h4a3;
			{8'd64, 8'd41}: color_data = 12'h4a3;
			{8'd64, 8'd42}: color_data = 12'h4b3;
			{8'd64, 8'd43}: color_data = 12'h4b3;
			{8'd64, 8'd44}: color_data = 12'h120;
			{8'd64, 8'd45}: color_data = 12'h000;
			{8'd64, 8'd46}: color_data = 12'h000;
			{8'd64, 8'd47}: color_data = 12'h000;
			{8'd64, 8'd48}: color_data = 12'h000;
			{8'd64, 8'd49}: color_data = 12'h000;
			{8'd64, 8'd50}: color_data = 12'h000;
			{8'd64, 8'd51}: color_data = 12'h000;
			{8'd64, 8'd52}: color_data = 12'h000;
			{8'd64, 8'd53}: color_data = 12'h382;
			{8'd64, 8'd54}: color_data = 12'h4b3;
			{8'd64, 8'd55}: color_data = 12'h4a3;
			{8'd64, 8'd56}: color_data = 12'h4a3;
			{8'd64, 8'd57}: color_data = 12'h4a3;
			{8'd64, 8'd58}: color_data = 12'h4a3;
			{8'd64, 8'd59}: color_data = 12'h4b3;
			{8'd64, 8'd60}: color_data = 12'h392;
			{8'd64, 8'd61}: color_data = 12'h000;
			{8'd64, 8'd62}: color_data = 12'h000;
			{8'd64, 8'd63}: color_data = 12'h000;
			{8'd64, 8'd64}: color_data = 12'h000;
			{8'd64, 8'd65}: color_data = 12'h000;
			{8'd64, 8'd66}: color_data = 12'h000;
			{8'd64, 8'd67}: color_data = 12'h000;
			{8'd64, 8'd100}: color_data = 12'he00;
			{8'd64, 8'd101}: color_data = 12'hf01;
			{8'd64, 8'd102}: color_data = 12'he00;
			{8'd64, 8'd103}: color_data = 12'he00;
			{8'd64, 8'd104}: color_data = 12'he00;
			{8'd64, 8'd105}: color_data = 12'he00;
			{8'd64, 8'd106}: color_data = 12'hc00;
			{8'd64, 8'd117}: color_data = 12'he00;
			{8'd64, 8'd118}: color_data = 12'he00;
			{8'd64, 8'd119}: color_data = 12'he00;
			{8'd64, 8'd120}: color_data = 12'he01;
			{8'd64, 8'd121}: color_data = 12'hf00;
			{8'd64, 8'd138}: color_data = 12'he00;
			{8'd64, 8'd139}: color_data = 12'he00;
			{8'd64, 8'd140}: color_data = 12'he00;
			{8'd64, 8'd141}: color_data = 12'he00;
			{8'd64, 8'd142}: color_data = 12'he00;
			{8'd64, 8'd143}: color_data = 12'he01;
			{8'd64, 8'd144}: color_data = 12'he00;
			{8'd65, 8'd4}: color_data = 12'h000;
			{8'd65, 8'd5}: color_data = 12'h000;
			{8'd65, 8'd6}: color_data = 12'h000;
			{8'd65, 8'd7}: color_data = 12'h000;
			{8'd65, 8'd8}: color_data = 12'h000;
			{8'd65, 8'd9}: color_data = 12'h000;
			{8'd65, 8'd10}: color_data = 12'h000;
			{8'd65, 8'd11}: color_data = 12'h000;
			{8'd65, 8'd12}: color_data = 12'h000;
			{8'd65, 8'd13}: color_data = 12'h000;
			{8'd65, 8'd14}: color_data = 12'h000;
			{8'd65, 8'd15}: color_data = 12'h000;
			{8'd65, 8'd16}: color_data = 12'h000;
			{8'd65, 8'd17}: color_data = 12'h000;
			{8'd65, 8'd18}: color_data = 12'h000;
			{8'd65, 8'd19}: color_data = 12'h000;
			{8'd65, 8'd20}: color_data = 12'h000;
			{8'd65, 8'd21}: color_data = 12'h000;
			{8'd65, 8'd22}: color_data = 12'h970;
			{8'd65, 8'd23}: color_data = 12'hfd0;
			{8'd65, 8'd24}: color_data = 12'hfc0;
			{8'd65, 8'd25}: color_data = 12'hfc0;
			{8'd65, 8'd26}: color_data = 12'hfc0;
			{8'd65, 8'd27}: color_data = 12'hfc0;
			{8'd65, 8'd28}: color_data = 12'hfd0;
			{8'd65, 8'd29}: color_data = 12'hfc0;
			{8'd65, 8'd30}: color_data = 12'h220;
			{8'd65, 8'd31}: color_data = 12'h000;
			{8'd65, 8'd32}: color_data = 12'h000;
			{8'd65, 8'd33}: color_data = 12'h000;
			{8'd65, 8'd34}: color_data = 12'h000;
			{8'd65, 8'd35}: color_data = 12'h272;
			{8'd65, 8'd36}: color_data = 12'h4b3;
			{8'd65, 8'd37}: color_data = 12'h4a3;
			{8'd65, 8'd38}: color_data = 12'h4a3;
			{8'd65, 8'd39}: color_data = 12'h4a3;
			{8'd65, 8'd40}: color_data = 12'h4a3;
			{8'd65, 8'd41}: color_data = 12'h4a3;
			{8'd65, 8'd42}: color_data = 12'h4a3;
			{8'd65, 8'd43}: color_data = 12'h4b3;
			{8'd65, 8'd44}: color_data = 12'h131;
			{8'd65, 8'd45}: color_data = 12'h000;
			{8'd65, 8'd46}: color_data = 12'h000;
			{8'd65, 8'd47}: color_data = 12'h000;
			{8'd65, 8'd48}: color_data = 12'h000;
			{8'd65, 8'd49}: color_data = 12'h000;
			{8'd65, 8'd50}: color_data = 12'h000;
			{8'd65, 8'd51}: color_data = 12'h000;
			{8'd65, 8'd52}: color_data = 12'h000;
			{8'd65, 8'd53}: color_data = 12'h382;
			{8'd65, 8'd54}: color_data = 12'h4b3;
			{8'd65, 8'd55}: color_data = 12'h4a3;
			{8'd65, 8'd56}: color_data = 12'h4a3;
			{8'd65, 8'd57}: color_data = 12'h4a3;
			{8'd65, 8'd58}: color_data = 12'h4a3;
			{8'd65, 8'd59}: color_data = 12'h4b3;
			{8'd65, 8'd60}: color_data = 12'h382;
			{8'd65, 8'd61}: color_data = 12'h000;
			{8'd65, 8'd62}: color_data = 12'h000;
			{8'd65, 8'd63}: color_data = 12'h000;
			{8'd65, 8'd64}: color_data = 12'h000;
			{8'd65, 8'd65}: color_data = 12'h000;
			{8'd65, 8'd66}: color_data = 12'h000;
			{8'd65, 8'd67}: color_data = 12'h000;
			{8'd65, 8'd100}: color_data = 12'he00;
			{8'd65, 8'd101}: color_data = 12'hf01;
			{8'd65, 8'd102}: color_data = 12'he00;
			{8'd65, 8'd103}: color_data = 12'he00;
			{8'd65, 8'd104}: color_data = 12'he00;
			{8'd65, 8'd105}: color_data = 12'he00;
			{8'd65, 8'd106}: color_data = 12'hc00;
			{8'd65, 8'd117}: color_data = 12'he00;
			{8'd65, 8'd118}: color_data = 12'he00;
			{8'd65, 8'd119}: color_data = 12'hf01;
			{8'd65, 8'd120}: color_data = 12'he00;
			{8'd65, 8'd121}: color_data = 12'he00;
			{8'd65, 8'd122}: color_data = 12'he00;
			{8'd65, 8'd123}: color_data = 12'he00;
			{8'd65, 8'd138}: color_data = 12'he00;
			{8'd65, 8'd139}: color_data = 12'he00;
			{8'd65, 8'd140}: color_data = 12'he00;
			{8'd65, 8'd141}: color_data = 12'he00;
			{8'd65, 8'd142}: color_data = 12'he00;
			{8'd65, 8'd143}: color_data = 12'he01;
			{8'd65, 8'd144}: color_data = 12'he00;
			{8'd66, 8'd4}: color_data = 12'h000;
			{8'd66, 8'd5}: color_data = 12'h000;
			{8'd66, 8'd6}: color_data = 12'h000;
			{8'd66, 8'd7}: color_data = 12'h000;
			{8'd66, 8'd8}: color_data = 12'h000;
			{8'd66, 8'd9}: color_data = 12'h000;
			{8'd66, 8'd10}: color_data = 12'h000;
			{8'd66, 8'd11}: color_data = 12'h000;
			{8'd66, 8'd12}: color_data = 12'h000;
			{8'd66, 8'd13}: color_data = 12'h000;
			{8'd66, 8'd14}: color_data = 12'h000;
			{8'd66, 8'd15}: color_data = 12'h000;
			{8'd66, 8'd16}: color_data = 12'h000;
			{8'd66, 8'd17}: color_data = 12'h000;
			{8'd66, 8'd18}: color_data = 12'h000;
			{8'd66, 8'd19}: color_data = 12'h000;
			{8'd66, 8'd20}: color_data = 12'h000;
			{8'd66, 8'd21}: color_data = 12'h000;
			{8'd66, 8'd22}: color_data = 12'ha80;
			{8'd66, 8'd23}: color_data = 12'hfd0;
			{8'd66, 8'd24}: color_data = 12'hfc0;
			{8'd66, 8'd25}: color_data = 12'hfc0;
			{8'd66, 8'd26}: color_data = 12'hfc0;
			{8'd66, 8'd27}: color_data = 12'hfc0;
			{8'd66, 8'd28}: color_data = 12'hfd0;
			{8'd66, 8'd29}: color_data = 12'hfc0;
			{8'd66, 8'd30}: color_data = 12'h220;
			{8'd66, 8'd31}: color_data = 12'h000;
			{8'd66, 8'd32}: color_data = 12'h000;
			{8'd66, 8'd33}: color_data = 12'h000;
			{8'd66, 8'd34}: color_data = 12'h000;
			{8'd66, 8'd35}: color_data = 12'h251;
			{8'd66, 8'd36}: color_data = 12'h4b3;
			{8'd66, 8'd37}: color_data = 12'h4a3;
			{8'd66, 8'd38}: color_data = 12'h4a3;
			{8'd66, 8'd39}: color_data = 12'h4a3;
			{8'd66, 8'd40}: color_data = 12'h4a3;
			{8'd66, 8'd41}: color_data = 12'h4a3;
			{8'd66, 8'd42}: color_data = 12'h4a3;
			{8'd66, 8'd43}: color_data = 12'h4b3;
			{8'd66, 8'd44}: color_data = 12'h272;
			{8'd66, 8'd45}: color_data = 12'h131;
			{8'd66, 8'd46}: color_data = 12'h010;
			{8'd66, 8'd47}: color_data = 12'h000;
			{8'd66, 8'd48}: color_data = 12'h000;
			{8'd66, 8'd49}: color_data = 12'h000;
			{8'd66, 8'd50}: color_data = 12'h000;
			{8'd66, 8'd51}: color_data = 12'h000;
			{8'd66, 8'd52}: color_data = 12'h000;
			{8'd66, 8'd53}: color_data = 12'h372;
			{8'd66, 8'd54}: color_data = 12'h4b3;
			{8'd66, 8'd55}: color_data = 12'h4a3;
			{8'd66, 8'd56}: color_data = 12'h4a3;
			{8'd66, 8'd57}: color_data = 12'h4a3;
			{8'd66, 8'd58}: color_data = 12'h4a3;
			{8'd66, 8'd59}: color_data = 12'h4b3;
			{8'd66, 8'd60}: color_data = 12'h262;
			{8'd66, 8'd61}: color_data = 12'h000;
			{8'd66, 8'd62}: color_data = 12'h000;
			{8'd66, 8'd63}: color_data = 12'h000;
			{8'd66, 8'd64}: color_data = 12'h000;
			{8'd66, 8'd65}: color_data = 12'h000;
			{8'd66, 8'd66}: color_data = 12'h000;
			{8'd66, 8'd67}: color_data = 12'h000;
			{8'd66, 8'd100}: color_data = 12'he00;
			{8'd66, 8'd101}: color_data = 12'hf01;
			{8'd66, 8'd102}: color_data = 12'he00;
			{8'd66, 8'd103}: color_data = 12'he00;
			{8'd66, 8'd104}: color_data = 12'he00;
			{8'd66, 8'd105}: color_data = 12'he00;
			{8'd66, 8'd106}: color_data = 12'hc00;
			{8'd66, 8'd117}: color_data = 12'he00;
			{8'd66, 8'd118}: color_data = 12'he00;
			{8'd66, 8'd119}: color_data = 12'he00;
			{8'd66, 8'd120}: color_data = 12'he00;
			{8'd66, 8'd121}: color_data = 12'he00;
			{8'd66, 8'd122}: color_data = 12'he01;
			{8'd66, 8'd123}: color_data = 12'he00;
			{8'd66, 8'd124}: color_data = 12'he00;
			{8'd66, 8'd125}: color_data = 12'he01;
			{8'd66, 8'd138}: color_data = 12'he00;
			{8'd66, 8'd139}: color_data = 12'he00;
			{8'd66, 8'd140}: color_data = 12'he00;
			{8'd66, 8'd141}: color_data = 12'he00;
			{8'd66, 8'd142}: color_data = 12'he00;
			{8'd66, 8'd143}: color_data = 12'he01;
			{8'd66, 8'd144}: color_data = 12'he00;
			{8'd67, 8'd6}: color_data = 12'h000;
			{8'd67, 8'd7}: color_data = 12'h000;
			{8'd67, 8'd8}: color_data = 12'h000;
			{8'd67, 8'd9}: color_data = 12'h000;
			{8'd67, 8'd10}: color_data = 12'h000;
			{8'd67, 8'd11}: color_data = 12'h000;
			{8'd67, 8'd12}: color_data = 12'h000;
			{8'd67, 8'd13}: color_data = 12'h000;
			{8'd67, 8'd14}: color_data = 12'h000;
			{8'd67, 8'd15}: color_data = 12'h000;
			{8'd67, 8'd16}: color_data = 12'h000;
			{8'd67, 8'd17}: color_data = 12'h000;
			{8'd67, 8'd18}: color_data = 12'h000;
			{8'd67, 8'd19}: color_data = 12'h000;
			{8'd67, 8'd20}: color_data = 12'h000;
			{8'd67, 8'd21}: color_data = 12'h000;
			{8'd67, 8'd22}: color_data = 12'hb90;
			{8'd67, 8'd23}: color_data = 12'hfd0;
			{8'd67, 8'd24}: color_data = 12'hfc0;
			{8'd67, 8'd25}: color_data = 12'hfc0;
			{8'd67, 8'd26}: color_data = 12'hfc0;
			{8'd67, 8'd27}: color_data = 12'hfc0;
			{8'd67, 8'd28}: color_data = 12'hfd0;
			{8'd67, 8'd29}: color_data = 12'hfc0;
			{8'd67, 8'd30}: color_data = 12'h320;
			{8'd67, 8'd31}: color_data = 12'h000;
			{8'd67, 8'd32}: color_data = 12'h000;
			{8'd67, 8'd33}: color_data = 12'h000;
			{8'd67, 8'd34}: color_data = 12'h000;
			{8'd67, 8'd35}: color_data = 12'h141;
			{8'd67, 8'd36}: color_data = 12'h4b3;
			{8'd67, 8'd37}: color_data = 12'h4a3;
			{8'd67, 8'd38}: color_data = 12'h4a3;
			{8'd67, 8'd39}: color_data = 12'h4a3;
			{8'd67, 8'd40}: color_data = 12'h4a3;
			{8'd67, 8'd41}: color_data = 12'h4a3;
			{8'd67, 8'd42}: color_data = 12'h4a3;
			{8'd67, 8'd43}: color_data = 12'h4a3;
			{8'd67, 8'd44}: color_data = 12'h4b3;
			{8'd67, 8'd45}: color_data = 12'h4b3;
			{8'd67, 8'd46}: color_data = 12'h4a3;
			{8'd67, 8'd47}: color_data = 12'h392;
			{8'd67, 8'd48}: color_data = 12'h272;
			{8'd67, 8'd49}: color_data = 12'h251;
			{8'd67, 8'd50}: color_data = 12'h130;
			{8'd67, 8'd51}: color_data = 12'h010;
			{8'd67, 8'd52}: color_data = 12'h000;
			{8'd67, 8'd53}: color_data = 12'h272;
			{8'd67, 8'd54}: color_data = 12'h4b3;
			{8'd67, 8'd55}: color_data = 12'h4a3;
			{8'd67, 8'd56}: color_data = 12'h4a3;
			{8'd67, 8'd57}: color_data = 12'h4a3;
			{8'd67, 8'd58}: color_data = 12'h4a3;
			{8'd67, 8'd59}: color_data = 12'h4b3;
			{8'd67, 8'd60}: color_data = 12'h151;
			{8'd67, 8'd61}: color_data = 12'h000;
			{8'd67, 8'd62}: color_data = 12'h000;
			{8'd67, 8'd63}: color_data = 12'h000;
			{8'd67, 8'd64}: color_data = 12'h000;
			{8'd67, 8'd65}: color_data = 12'h000;
			{8'd67, 8'd66}: color_data = 12'h000;
			{8'd67, 8'd67}: color_data = 12'h000;
			{8'd67, 8'd68}: color_data = 12'h000;
			{8'd67, 8'd69}: color_data = 12'h000;
			{8'd67, 8'd100}: color_data = 12'he00;
			{8'd67, 8'd101}: color_data = 12'hf01;
			{8'd67, 8'd102}: color_data = 12'he00;
			{8'd67, 8'd103}: color_data = 12'he00;
			{8'd67, 8'd104}: color_data = 12'he00;
			{8'd67, 8'd105}: color_data = 12'he00;
			{8'd67, 8'd106}: color_data = 12'hc00;
			{8'd67, 8'd117}: color_data = 12'he00;
			{8'd67, 8'd118}: color_data = 12'he00;
			{8'd67, 8'd119}: color_data = 12'he00;
			{8'd67, 8'd120}: color_data = 12'he00;
			{8'd67, 8'd121}: color_data = 12'he00;
			{8'd67, 8'd122}: color_data = 12'he00;
			{8'd67, 8'd123}: color_data = 12'he00;
			{8'd67, 8'd124}: color_data = 12'he01;
			{8'd67, 8'd125}: color_data = 12'he00;
			{8'd67, 8'd126}: color_data = 12'he00;
			{8'd67, 8'd127}: color_data = 12'he01;
			{8'd67, 8'd128}: color_data = 12'he01;
			{8'd67, 8'd138}: color_data = 12'he00;
			{8'd67, 8'd139}: color_data = 12'he00;
			{8'd67, 8'd140}: color_data = 12'he00;
			{8'd67, 8'd141}: color_data = 12'he00;
			{8'd67, 8'd142}: color_data = 12'he00;
			{8'd67, 8'd143}: color_data = 12'he01;
			{8'd67, 8'd144}: color_data = 12'he00;
			{8'd68, 8'd7}: color_data = 12'h000;
			{8'd68, 8'd8}: color_data = 12'h000;
			{8'd68, 8'd9}: color_data = 12'h540;
			{8'd68, 8'd10}: color_data = 12'heb0;
			{8'd68, 8'd11}: color_data = 12'hda0;
			{8'd68, 8'd12}: color_data = 12'hca0;
			{8'd68, 8'd13}: color_data = 12'hca0;
			{8'd68, 8'd14}: color_data = 12'hb90;
			{8'd68, 8'd15}: color_data = 12'ha80;
			{8'd68, 8'd16}: color_data = 12'ha80;
			{8'd68, 8'd17}: color_data = 12'h970;
			{8'd68, 8'd18}: color_data = 12'h870;
			{8'd68, 8'd19}: color_data = 12'h860;
			{8'd68, 8'd20}: color_data = 12'h760;
			{8'd68, 8'd21}: color_data = 12'h650;
			{8'd68, 8'd22}: color_data = 12'hdb0;
			{8'd68, 8'd23}: color_data = 12'hfd0;
			{8'd68, 8'd24}: color_data = 12'hfc0;
			{8'd68, 8'd25}: color_data = 12'hfc0;
			{8'd68, 8'd26}: color_data = 12'hfc0;
			{8'd68, 8'd27}: color_data = 12'hfc0;
			{8'd68, 8'd28}: color_data = 12'hfd0;
			{8'd68, 8'd29}: color_data = 12'hfd0;
			{8'd68, 8'd30}: color_data = 12'h320;
			{8'd68, 8'd31}: color_data = 12'h000;
			{8'd68, 8'd32}: color_data = 12'h000;
			{8'd68, 8'd33}: color_data = 12'h000;
			{8'd68, 8'd34}: color_data = 12'h000;
			{8'd68, 8'd35}: color_data = 12'h131;
			{8'd68, 8'd36}: color_data = 12'h4b3;
			{8'd68, 8'd37}: color_data = 12'h4a3;
			{8'd68, 8'd38}: color_data = 12'h4a3;
			{8'd68, 8'd39}: color_data = 12'h4a3;
			{8'd68, 8'd40}: color_data = 12'h4a3;
			{8'd68, 8'd41}: color_data = 12'h4a3;
			{8'd68, 8'd42}: color_data = 12'h4a3;
			{8'd68, 8'd43}: color_data = 12'h4a3;
			{8'd68, 8'd44}: color_data = 12'h4a3;
			{8'd68, 8'd45}: color_data = 12'h4a3;
			{8'd68, 8'd46}: color_data = 12'h4b3;
			{8'd68, 8'd47}: color_data = 12'h4b3;
			{8'd68, 8'd48}: color_data = 12'h4b3;
			{8'd68, 8'd49}: color_data = 12'h4b3;
			{8'd68, 8'd50}: color_data = 12'h4b3;
			{8'd68, 8'd51}: color_data = 12'h4a3;
			{8'd68, 8'd52}: color_data = 12'h382;
			{8'd68, 8'd53}: color_data = 12'h392;
			{8'd68, 8'd54}: color_data = 12'h4b3;
			{8'd68, 8'd55}: color_data = 12'h4a3;
			{8'd68, 8'd56}: color_data = 12'h4a3;
			{8'd68, 8'd57}: color_data = 12'h4a3;
			{8'd68, 8'd58}: color_data = 12'h4a3;
			{8'd68, 8'd59}: color_data = 12'h4b3;
			{8'd68, 8'd60}: color_data = 12'h131;
			{8'd68, 8'd61}: color_data = 12'h000;
			{8'd68, 8'd62}: color_data = 12'h000;
			{8'd68, 8'd63}: color_data = 12'h000;
			{8'd68, 8'd64}: color_data = 12'h000;
			{8'd68, 8'd65}: color_data = 12'h000;
			{8'd68, 8'd66}: color_data = 12'h000;
			{8'd68, 8'd67}: color_data = 12'h000;
			{8'd68, 8'd68}: color_data = 12'h000;
			{8'd68, 8'd69}: color_data = 12'h000;
			{8'd68, 8'd70}: color_data = 12'h000;
			{8'd68, 8'd71}: color_data = 12'h000;
			{8'd68, 8'd72}: color_data = 12'h000;
			{8'd68, 8'd73}: color_data = 12'h000;
			{8'd68, 8'd74}: color_data = 12'h000;
			{8'd68, 8'd100}: color_data = 12'he00;
			{8'd68, 8'd101}: color_data = 12'hf01;
			{8'd68, 8'd102}: color_data = 12'he00;
			{8'd68, 8'd103}: color_data = 12'he00;
			{8'd68, 8'd104}: color_data = 12'he00;
			{8'd68, 8'd105}: color_data = 12'he00;
			{8'd68, 8'd106}: color_data = 12'hc00;
			{8'd68, 8'd117}: color_data = 12'he00;
			{8'd68, 8'd118}: color_data = 12'he00;
			{8'd68, 8'd119}: color_data = 12'he00;
			{8'd68, 8'd120}: color_data = 12'he00;
			{8'd68, 8'd121}: color_data = 12'he00;
			{8'd68, 8'd122}: color_data = 12'he00;
			{8'd68, 8'd123}: color_data = 12'he00;
			{8'd68, 8'd124}: color_data = 12'he00;
			{8'd68, 8'd125}: color_data = 12'he00;
			{8'd68, 8'd126}: color_data = 12'he01;
			{8'd68, 8'd127}: color_data = 12'he00;
			{8'd68, 8'd128}: color_data = 12'he00;
			{8'd68, 8'd129}: color_data = 12'he00;
			{8'd68, 8'd130}: color_data = 12'he01;
			{8'd68, 8'd138}: color_data = 12'he00;
			{8'd68, 8'd139}: color_data = 12'he00;
			{8'd68, 8'd140}: color_data = 12'he00;
			{8'd68, 8'd141}: color_data = 12'he00;
			{8'd68, 8'd142}: color_data = 12'he00;
			{8'd68, 8'd143}: color_data = 12'he01;
			{8'd68, 8'd144}: color_data = 12'he00;
			{8'd69, 8'd7}: color_data = 12'h000;
			{8'd69, 8'd8}: color_data = 12'h000;
			{8'd69, 8'd9}: color_data = 12'h540;
			{8'd69, 8'd10}: color_data = 12'hfd0;
			{8'd69, 8'd11}: color_data = 12'hfd0;
			{8'd69, 8'd12}: color_data = 12'hfd0;
			{8'd69, 8'd13}: color_data = 12'hfd0;
			{8'd69, 8'd14}: color_data = 12'hfd0;
			{8'd69, 8'd15}: color_data = 12'hfd0;
			{8'd69, 8'd16}: color_data = 12'hfd0;
			{8'd69, 8'd17}: color_data = 12'hfd0;
			{8'd69, 8'd18}: color_data = 12'hfd0;
			{8'd69, 8'd19}: color_data = 12'hfd0;
			{8'd69, 8'd20}: color_data = 12'hfd0;
			{8'd69, 8'd21}: color_data = 12'hfd0;
			{8'd69, 8'd22}: color_data = 12'hfd0;
			{8'd69, 8'd23}: color_data = 12'hfc0;
			{8'd69, 8'd24}: color_data = 12'hfc0;
			{8'd69, 8'd25}: color_data = 12'hfc0;
			{8'd69, 8'd26}: color_data = 12'hfc0;
			{8'd69, 8'd27}: color_data = 12'hfc0;
			{8'd69, 8'd28}: color_data = 12'hfd0;
			{8'd69, 8'd29}: color_data = 12'hfd0;
			{8'd69, 8'd30}: color_data = 12'h330;
			{8'd69, 8'd31}: color_data = 12'h000;
			{8'd69, 8'd32}: color_data = 12'h000;
			{8'd69, 8'd33}: color_data = 12'h000;
			{8'd69, 8'd34}: color_data = 12'h000;
			{8'd69, 8'd35}: color_data = 12'h120;
			{8'd69, 8'd36}: color_data = 12'h4b3;
			{8'd69, 8'd37}: color_data = 12'h4a3;
			{8'd69, 8'd38}: color_data = 12'h4a3;
			{8'd69, 8'd39}: color_data = 12'h4a3;
			{8'd69, 8'd40}: color_data = 12'h4a3;
			{8'd69, 8'd41}: color_data = 12'h4a3;
			{8'd69, 8'd42}: color_data = 12'h4a3;
			{8'd69, 8'd43}: color_data = 12'h4a3;
			{8'd69, 8'd44}: color_data = 12'h4a3;
			{8'd69, 8'd45}: color_data = 12'h4a3;
			{8'd69, 8'd46}: color_data = 12'h4a3;
			{8'd69, 8'd47}: color_data = 12'h4a3;
			{8'd69, 8'd48}: color_data = 12'h4a3;
			{8'd69, 8'd49}: color_data = 12'h4a3;
			{8'd69, 8'd50}: color_data = 12'h4a3;
			{8'd69, 8'd51}: color_data = 12'h4b3;
			{8'd69, 8'd52}: color_data = 12'h4b3;
			{8'd69, 8'd53}: color_data = 12'h4b3;
			{8'd69, 8'd54}: color_data = 12'h4a3;
			{8'd69, 8'd55}: color_data = 12'h4a3;
			{8'd69, 8'd56}: color_data = 12'h4a3;
			{8'd69, 8'd57}: color_data = 12'h4a3;
			{8'd69, 8'd58}: color_data = 12'h4b3;
			{8'd69, 8'd59}: color_data = 12'h4a3;
			{8'd69, 8'd60}: color_data = 12'h131;
			{8'd69, 8'd61}: color_data = 12'h000;
			{8'd69, 8'd62}: color_data = 12'h000;
			{8'd69, 8'd63}: color_data = 12'h000;
			{8'd69, 8'd64}: color_data = 12'h000;
			{8'd69, 8'd65}: color_data = 12'h000;
			{8'd69, 8'd66}: color_data = 12'h000;
			{8'd69, 8'd67}: color_data = 12'h000;
			{8'd69, 8'd68}: color_data = 12'h000;
			{8'd69, 8'd69}: color_data = 12'h000;
			{8'd69, 8'd70}: color_data = 12'h000;
			{8'd69, 8'd71}: color_data = 12'h000;
			{8'd69, 8'd72}: color_data = 12'h000;
			{8'd69, 8'd73}: color_data = 12'h000;
			{8'd69, 8'd74}: color_data = 12'h000;
			{8'd69, 8'd75}: color_data = 12'h000;
			{8'd69, 8'd100}: color_data = 12'he00;
			{8'd69, 8'd101}: color_data = 12'hf01;
			{8'd69, 8'd102}: color_data = 12'he00;
			{8'd69, 8'd103}: color_data = 12'he00;
			{8'd69, 8'd104}: color_data = 12'he00;
			{8'd69, 8'd105}: color_data = 12'he00;
			{8'd69, 8'd106}: color_data = 12'hc00;
			{8'd69, 8'd117}: color_data = 12'he01;
			{8'd69, 8'd118}: color_data = 12'he00;
			{8'd69, 8'd119}: color_data = 12'hf01;
			{8'd69, 8'd120}: color_data = 12'he00;
			{8'd69, 8'd121}: color_data = 12'he00;
			{8'd69, 8'd122}: color_data = 12'he00;
			{8'd69, 8'd123}: color_data = 12'he00;
			{8'd69, 8'd124}: color_data = 12'he00;
			{8'd69, 8'd125}: color_data = 12'he00;
			{8'd69, 8'd126}: color_data = 12'he00;
			{8'd69, 8'd127}: color_data = 12'he00;
			{8'd69, 8'd128}: color_data = 12'he00;
			{8'd69, 8'd129}: color_data = 12'he01;
			{8'd69, 8'd130}: color_data = 12'he00;
			{8'd69, 8'd131}: color_data = 12'he00;
			{8'd69, 8'd132}: color_data = 12'he01;
			{8'd69, 8'd133}: color_data = 12'ha00;
			{8'd69, 8'd138}: color_data = 12'he00;
			{8'd69, 8'd139}: color_data = 12'he00;
			{8'd69, 8'd140}: color_data = 12'he00;
			{8'd69, 8'd141}: color_data = 12'he00;
			{8'd69, 8'd142}: color_data = 12'he00;
			{8'd69, 8'd143}: color_data = 12'he01;
			{8'd69, 8'd144}: color_data = 12'he00;
			{8'd70, 8'd7}: color_data = 12'h000;
			{8'd70, 8'd8}: color_data = 12'h000;
			{8'd70, 8'd9}: color_data = 12'h320;
			{8'd70, 8'd10}: color_data = 12'hfc0;
			{8'd70, 8'd11}: color_data = 12'hfd0;
			{8'd70, 8'd12}: color_data = 12'hfc0;
			{8'd70, 8'd13}: color_data = 12'hfc0;
			{8'd70, 8'd14}: color_data = 12'hfc0;
			{8'd70, 8'd15}: color_data = 12'hfc0;
			{8'd70, 8'd16}: color_data = 12'hfc0;
			{8'd70, 8'd17}: color_data = 12'hfc0;
			{8'd70, 8'd18}: color_data = 12'hfc0;
			{8'd70, 8'd19}: color_data = 12'hfc0;
			{8'd70, 8'd20}: color_data = 12'hfc0;
			{8'd70, 8'd21}: color_data = 12'hfc0;
			{8'd70, 8'd22}: color_data = 12'hfc0;
			{8'd70, 8'd23}: color_data = 12'hfc0;
			{8'd70, 8'd24}: color_data = 12'hfc0;
			{8'd70, 8'd25}: color_data = 12'hfc0;
			{8'd70, 8'd26}: color_data = 12'hfc0;
			{8'd70, 8'd27}: color_data = 12'hfc0;
			{8'd70, 8'd28}: color_data = 12'hfd0;
			{8'd70, 8'd29}: color_data = 12'hfd0;
			{8'd70, 8'd30}: color_data = 12'h330;
			{8'd70, 8'd31}: color_data = 12'h000;
			{8'd70, 8'd32}: color_data = 12'h000;
			{8'd70, 8'd33}: color_data = 12'h000;
			{8'd70, 8'd34}: color_data = 12'h000;
			{8'd70, 8'd35}: color_data = 12'h010;
			{8'd70, 8'd36}: color_data = 12'h4a3;
			{8'd70, 8'd37}: color_data = 12'h4b3;
			{8'd70, 8'd38}: color_data = 12'h4a3;
			{8'd70, 8'd39}: color_data = 12'h4a3;
			{8'd70, 8'd40}: color_data = 12'h4a3;
			{8'd70, 8'd41}: color_data = 12'h4a3;
			{8'd70, 8'd42}: color_data = 12'h4a3;
			{8'd70, 8'd43}: color_data = 12'h4a3;
			{8'd70, 8'd44}: color_data = 12'h4a3;
			{8'd70, 8'd45}: color_data = 12'h4a3;
			{8'd70, 8'd46}: color_data = 12'h4a3;
			{8'd70, 8'd47}: color_data = 12'h4a3;
			{8'd70, 8'd48}: color_data = 12'h4a3;
			{8'd70, 8'd49}: color_data = 12'h4a3;
			{8'd70, 8'd50}: color_data = 12'h4a3;
			{8'd70, 8'd51}: color_data = 12'h4a3;
			{8'd70, 8'd52}: color_data = 12'h4a3;
			{8'd70, 8'd53}: color_data = 12'h4a3;
			{8'd70, 8'd54}: color_data = 12'h4a3;
			{8'd70, 8'd55}: color_data = 12'h4a3;
			{8'd70, 8'd56}: color_data = 12'h4a3;
			{8'd70, 8'd57}: color_data = 12'h4a3;
			{8'd70, 8'd58}: color_data = 12'h4a3;
			{8'd70, 8'd59}: color_data = 12'h4a3;
			{8'd70, 8'd60}: color_data = 12'h4a3;
			{8'd70, 8'd61}: color_data = 12'h393;
			{8'd70, 8'd62}: color_data = 12'h382;
			{8'd70, 8'd63}: color_data = 12'h261;
			{8'd70, 8'd64}: color_data = 12'h141;
			{8'd70, 8'd65}: color_data = 12'h020;
			{8'd70, 8'd66}: color_data = 12'h000;
			{8'd70, 8'd67}: color_data = 12'h000;
			{8'd70, 8'd68}: color_data = 12'h000;
			{8'd70, 8'd69}: color_data = 12'h000;
			{8'd70, 8'd70}: color_data = 12'h000;
			{8'd70, 8'd71}: color_data = 12'h000;
			{8'd70, 8'd72}: color_data = 12'h000;
			{8'd70, 8'd73}: color_data = 12'h000;
			{8'd70, 8'd74}: color_data = 12'h000;
			{8'd70, 8'd75}: color_data = 12'h000;
			{8'd70, 8'd100}: color_data = 12'he00;
			{8'd70, 8'd101}: color_data = 12'hf01;
			{8'd70, 8'd102}: color_data = 12'he00;
			{8'd70, 8'd103}: color_data = 12'he00;
			{8'd70, 8'd104}: color_data = 12'he00;
			{8'd70, 8'd105}: color_data = 12'he00;
			{8'd70, 8'd106}: color_data = 12'hc00;
			{8'd70, 8'd117}: color_data = 12'hf00;
			{8'd70, 8'd118}: color_data = 12'he00;
			{8'd70, 8'd119}: color_data = 12'he00;
			{8'd70, 8'd120}: color_data = 12'he00;
			{8'd70, 8'd121}: color_data = 12'he00;
			{8'd70, 8'd122}: color_data = 12'he01;
			{8'd70, 8'd123}: color_data = 12'he00;
			{8'd70, 8'd124}: color_data = 12'he00;
			{8'd70, 8'd125}: color_data = 12'he00;
			{8'd70, 8'd126}: color_data = 12'he00;
			{8'd70, 8'd127}: color_data = 12'he00;
			{8'd70, 8'd128}: color_data = 12'he00;
			{8'd70, 8'd129}: color_data = 12'he00;
			{8'd70, 8'd130}: color_data = 12'he00;
			{8'd70, 8'd131}: color_data = 12'he01;
			{8'd70, 8'd132}: color_data = 12'he00;
			{8'd70, 8'd133}: color_data = 12'he00;
			{8'd70, 8'd138}: color_data = 12'he00;
			{8'd70, 8'd139}: color_data = 12'he00;
			{8'd70, 8'd140}: color_data = 12'he00;
			{8'd70, 8'd141}: color_data = 12'he00;
			{8'd70, 8'd142}: color_data = 12'he00;
			{8'd70, 8'd143}: color_data = 12'he01;
			{8'd70, 8'd144}: color_data = 12'he00;
			{8'd71, 8'd7}: color_data = 12'h000;
			{8'd71, 8'd8}: color_data = 12'h000;
			{8'd71, 8'd9}: color_data = 12'h110;
			{8'd71, 8'd10}: color_data = 12'hec0;
			{8'd71, 8'd11}: color_data = 12'hfd0;
			{8'd71, 8'd12}: color_data = 12'hfc0;
			{8'd71, 8'd13}: color_data = 12'hfc0;
			{8'd71, 8'd14}: color_data = 12'hfc0;
			{8'd71, 8'd15}: color_data = 12'hfc0;
			{8'd71, 8'd16}: color_data = 12'hfc0;
			{8'd71, 8'd17}: color_data = 12'hfc0;
			{8'd71, 8'd18}: color_data = 12'hfc0;
			{8'd71, 8'd19}: color_data = 12'hfc0;
			{8'd71, 8'd20}: color_data = 12'hfc0;
			{8'd71, 8'd21}: color_data = 12'hfc0;
			{8'd71, 8'd22}: color_data = 12'hfc0;
			{8'd71, 8'd23}: color_data = 12'hfc0;
			{8'd71, 8'd24}: color_data = 12'hfc0;
			{8'd71, 8'd25}: color_data = 12'hfc0;
			{8'd71, 8'd26}: color_data = 12'hfc0;
			{8'd71, 8'd27}: color_data = 12'hfd0;
			{8'd71, 8'd28}: color_data = 12'hfd0;
			{8'd71, 8'd29}: color_data = 12'ha80;
			{8'd71, 8'd30}: color_data = 12'h000;
			{8'd71, 8'd31}: color_data = 12'h000;
			{8'd71, 8'd32}: color_data = 12'h000;
			{8'd71, 8'd33}: color_data = 12'h000;
			{8'd71, 8'd34}: color_data = 12'h000;
			{8'd71, 8'd35}: color_data = 12'h000;
			{8'd71, 8'd36}: color_data = 12'h393;
			{8'd71, 8'd37}: color_data = 12'h4b3;
			{8'd71, 8'd38}: color_data = 12'h4b3;
			{8'd71, 8'd39}: color_data = 12'h4b3;
			{8'd71, 8'd40}: color_data = 12'h4a3;
			{8'd71, 8'd41}: color_data = 12'h4a3;
			{8'd71, 8'd42}: color_data = 12'h4a3;
			{8'd71, 8'd43}: color_data = 12'h4a3;
			{8'd71, 8'd44}: color_data = 12'h4a3;
			{8'd71, 8'd45}: color_data = 12'h4a3;
			{8'd71, 8'd46}: color_data = 12'h4a3;
			{8'd71, 8'd47}: color_data = 12'h4a3;
			{8'd71, 8'd48}: color_data = 12'h4a3;
			{8'd71, 8'd49}: color_data = 12'h4a3;
			{8'd71, 8'd50}: color_data = 12'h4a3;
			{8'd71, 8'd51}: color_data = 12'h4a3;
			{8'd71, 8'd52}: color_data = 12'h4a3;
			{8'd71, 8'd53}: color_data = 12'h4a3;
			{8'd71, 8'd54}: color_data = 12'h4a3;
			{8'd71, 8'd55}: color_data = 12'h4a3;
			{8'd71, 8'd56}: color_data = 12'h4a3;
			{8'd71, 8'd57}: color_data = 12'h4a3;
			{8'd71, 8'd58}: color_data = 12'h4a3;
			{8'd71, 8'd59}: color_data = 12'h4a3;
			{8'd71, 8'd60}: color_data = 12'h4b3;
			{8'd71, 8'd61}: color_data = 12'h4b3;
			{8'd71, 8'd62}: color_data = 12'h4b3;
			{8'd71, 8'd63}: color_data = 12'h4b3;
			{8'd71, 8'd64}: color_data = 12'h4b3;
			{8'd71, 8'd65}: color_data = 12'h4a3;
			{8'd71, 8'd66}: color_data = 12'h392;
			{8'd71, 8'd67}: color_data = 12'h272;
			{8'd71, 8'd68}: color_data = 12'h000;
			{8'd71, 8'd69}: color_data = 12'h000;
			{8'd71, 8'd70}: color_data = 12'h000;
			{8'd71, 8'd71}: color_data = 12'h000;
			{8'd71, 8'd72}: color_data = 12'h000;
			{8'd71, 8'd73}: color_data = 12'h000;
			{8'd71, 8'd74}: color_data = 12'h000;
			{8'd71, 8'd75}: color_data = 12'h000;
			{8'd71, 8'd100}: color_data = 12'he00;
			{8'd71, 8'd101}: color_data = 12'hf01;
			{8'd71, 8'd102}: color_data = 12'he00;
			{8'd71, 8'd103}: color_data = 12'he00;
			{8'd71, 8'd104}: color_data = 12'he00;
			{8'd71, 8'd105}: color_data = 12'he00;
			{8'd71, 8'd106}: color_data = 12'hc00;
			{8'd71, 8'd120}: color_data = 12'hf00;
			{8'd71, 8'd121}: color_data = 12'he00;
			{8'd71, 8'd122}: color_data = 12'he00;
			{8'd71, 8'd123}: color_data = 12'he00;
			{8'd71, 8'd124}: color_data = 12'he00;
			{8'd71, 8'd125}: color_data = 12'he00;
			{8'd71, 8'd126}: color_data = 12'he01;
			{8'd71, 8'd127}: color_data = 12'he00;
			{8'd71, 8'd128}: color_data = 12'he00;
			{8'd71, 8'd129}: color_data = 12'he00;
			{8'd71, 8'd130}: color_data = 12'he00;
			{8'd71, 8'd131}: color_data = 12'he00;
			{8'd71, 8'd132}: color_data = 12'hf01;
			{8'd71, 8'd133}: color_data = 12'he00;
			{8'd71, 8'd138}: color_data = 12'he00;
			{8'd71, 8'd139}: color_data = 12'he00;
			{8'd71, 8'd140}: color_data = 12'he00;
			{8'd71, 8'd141}: color_data = 12'he00;
			{8'd71, 8'd142}: color_data = 12'he00;
			{8'd71, 8'd143}: color_data = 12'he01;
			{8'd71, 8'd144}: color_data = 12'he00;
			{8'd72, 8'd7}: color_data = 12'h000;
			{8'd72, 8'd8}: color_data = 12'h000;
			{8'd72, 8'd9}: color_data = 12'h000;
			{8'd72, 8'd10}: color_data = 12'hdb0;
			{8'd72, 8'd11}: color_data = 12'hfd0;
			{8'd72, 8'd12}: color_data = 12'hfc0;
			{8'd72, 8'd13}: color_data = 12'hfc0;
			{8'd72, 8'd14}: color_data = 12'hfc0;
			{8'd72, 8'd15}: color_data = 12'hfc0;
			{8'd72, 8'd16}: color_data = 12'hfc0;
			{8'd72, 8'd17}: color_data = 12'hfc0;
			{8'd72, 8'd18}: color_data = 12'hfc0;
			{8'd72, 8'd19}: color_data = 12'hfc0;
			{8'd72, 8'd20}: color_data = 12'hfc0;
			{8'd72, 8'd21}: color_data = 12'hfc0;
			{8'd72, 8'd22}: color_data = 12'hfc0;
			{8'd72, 8'd23}: color_data = 12'hfc0;
			{8'd72, 8'd24}: color_data = 12'hfc0;
			{8'd72, 8'd25}: color_data = 12'hfc0;
			{8'd72, 8'd26}: color_data = 12'hfd0;
			{8'd72, 8'd27}: color_data = 12'hfd0;
			{8'd72, 8'd28}: color_data = 12'h970;
			{8'd72, 8'd29}: color_data = 12'h000;
			{8'd72, 8'd30}: color_data = 12'h000;
			{8'd72, 8'd31}: color_data = 12'h000;
			{8'd72, 8'd32}: color_data = 12'h000;
			{8'd72, 8'd33}: color_data = 12'h000;
			{8'd72, 8'd34}: color_data = 12'h000;
			{8'd72, 8'd35}: color_data = 12'h000;
			{8'd72, 8'd36}: color_data = 12'h010;
			{8'd72, 8'd37}: color_data = 12'h251;
			{8'd72, 8'd38}: color_data = 12'h392;
			{8'd72, 8'd39}: color_data = 12'h4b3;
			{8'd72, 8'd40}: color_data = 12'h4b3;
			{8'd72, 8'd41}: color_data = 12'h4b3;
			{8'd72, 8'd42}: color_data = 12'h4b3;
			{8'd72, 8'd43}: color_data = 12'h4a3;
			{8'd72, 8'd44}: color_data = 12'h4a3;
			{8'd72, 8'd45}: color_data = 12'h4a3;
			{8'd72, 8'd46}: color_data = 12'h4a3;
			{8'd72, 8'd47}: color_data = 12'h4a3;
			{8'd72, 8'd48}: color_data = 12'h4a3;
			{8'd72, 8'd49}: color_data = 12'h4a3;
			{8'd72, 8'd50}: color_data = 12'h4a3;
			{8'd72, 8'd51}: color_data = 12'h4a3;
			{8'd72, 8'd52}: color_data = 12'h4a3;
			{8'd72, 8'd53}: color_data = 12'h4a3;
			{8'd72, 8'd54}: color_data = 12'h4a3;
			{8'd72, 8'd55}: color_data = 12'h4a3;
			{8'd72, 8'd56}: color_data = 12'h4a3;
			{8'd72, 8'd57}: color_data = 12'h4a3;
			{8'd72, 8'd58}: color_data = 12'h4a3;
			{8'd72, 8'd59}: color_data = 12'h4a3;
			{8'd72, 8'd60}: color_data = 12'h4a3;
			{8'd72, 8'd61}: color_data = 12'h4a3;
			{8'd72, 8'd62}: color_data = 12'h4a3;
			{8'd72, 8'd63}: color_data = 12'h4a3;
			{8'd72, 8'd64}: color_data = 12'h4a3;
			{8'd72, 8'd65}: color_data = 12'h4b3;
			{8'd72, 8'd66}: color_data = 12'h4b3;
			{8'd72, 8'd67}: color_data = 12'h4a3;
			{8'd72, 8'd68}: color_data = 12'h000;
			{8'd72, 8'd69}: color_data = 12'h000;
			{8'd72, 8'd70}: color_data = 12'h000;
			{8'd72, 8'd71}: color_data = 12'h000;
			{8'd72, 8'd72}: color_data = 12'h000;
			{8'd72, 8'd73}: color_data = 12'h000;
			{8'd72, 8'd74}: color_data = 12'h000;
			{8'd72, 8'd100}: color_data = 12'he00;
			{8'd72, 8'd101}: color_data = 12'hf01;
			{8'd72, 8'd102}: color_data = 12'he00;
			{8'd72, 8'd103}: color_data = 12'he00;
			{8'd72, 8'd104}: color_data = 12'he00;
			{8'd72, 8'd105}: color_data = 12'he00;
			{8'd72, 8'd106}: color_data = 12'hc00;
			{8'd72, 8'd124}: color_data = 12'he00;
			{8'd72, 8'd125}: color_data = 12'he00;
			{8'd72, 8'd126}: color_data = 12'he00;
			{8'd72, 8'd127}: color_data = 12'he00;
			{8'd72, 8'd128}: color_data = 12'he00;
			{8'd72, 8'd129}: color_data = 12'he00;
			{8'd72, 8'd130}: color_data = 12'he00;
			{8'd72, 8'd131}: color_data = 12'he00;
			{8'd72, 8'd132}: color_data = 12'hf01;
			{8'd72, 8'd133}: color_data = 12'he00;
			{8'd72, 8'd138}: color_data = 12'he00;
			{8'd72, 8'd139}: color_data = 12'he00;
			{8'd72, 8'd140}: color_data = 12'he00;
			{8'd72, 8'd141}: color_data = 12'he00;
			{8'd72, 8'd142}: color_data = 12'he00;
			{8'd72, 8'd143}: color_data = 12'he01;
			{8'd72, 8'd144}: color_data = 12'he00;
			{8'd73, 8'd7}: color_data = 12'h000;
			{8'd73, 8'd8}: color_data = 12'h000;
			{8'd73, 8'd9}: color_data = 12'h000;
			{8'd73, 8'd10}: color_data = 12'hca0;
			{8'd73, 8'd11}: color_data = 12'hfd0;
			{8'd73, 8'd12}: color_data = 12'hfc0;
			{8'd73, 8'd13}: color_data = 12'hfc0;
			{8'd73, 8'd14}: color_data = 12'hfc0;
			{8'd73, 8'd15}: color_data = 12'hfc0;
			{8'd73, 8'd16}: color_data = 12'hfc0;
			{8'd73, 8'd17}: color_data = 12'hfc0;
			{8'd73, 8'd18}: color_data = 12'hfc0;
			{8'd73, 8'd19}: color_data = 12'hfc0;
			{8'd73, 8'd20}: color_data = 12'hfc0;
			{8'd73, 8'd21}: color_data = 12'hfc0;
			{8'd73, 8'd22}: color_data = 12'hfc0;
			{8'd73, 8'd23}: color_data = 12'hfc0;
			{8'd73, 8'd24}: color_data = 12'hfc0;
			{8'd73, 8'd25}: color_data = 12'hfd0;
			{8'd73, 8'd26}: color_data = 12'hfd0;
			{8'd73, 8'd27}: color_data = 12'h760;
			{8'd73, 8'd28}: color_data = 12'h000;
			{8'd73, 8'd29}: color_data = 12'h000;
			{8'd73, 8'd30}: color_data = 12'h000;
			{8'd73, 8'd31}: color_data = 12'h000;
			{8'd73, 8'd32}: color_data = 12'h000;
			{8'd73, 8'd33}: color_data = 12'h000;
			{8'd73, 8'd34}: color_data = 12'h000;
			{8'd73, 8'd35}: color_data = 12'h000;
			{8'd73, 8'd36}: color_data = 12'h000;
			{8'd73, 8'd37}: color_data = 12'h000;
			{8'd73, 8'd38}: color_data = 12'h000;
			{8'd73, 8'd39}: color_data = 12'h120;
			{8'd73, 8'd40}: color_data = 12'h261;
			{8'd73, 8'd41}: color_data = 12'h392;
			{8'd73, 8'd42}: color_data = 12'h4b3;
			{8'd73, 8'd43}: color_data = 12'h4b3;
			{8'd73, 8'd44}: color_data = 12'h4b3;
			{8'd73, 8'd45}: color_data = 12'h4a3;
			{8'd73, 8'd46}: color_data = 12'h4a3;
			{8'd73, 8'd47}: color_data = 12'h4a3;
			{8'd73, 8'd48}: color_data = 12'h4a3;
			{8'd73, 8'd49}: color_data = 12'h4a3;
			{8'd73, 8'd50}: color_data = 12'h4a3;
			{8'd73, 8'd51}: color_data = 12'h4a3;
			{8'd73, 8'd52}: color_data = 12'h4a3;
			{8'd73, 8'd53}: color_data = 12'h4a3;
			{8'd73, 8'd54}: color_data = 12'h4a3;
			{8'd73, 8'd55}: color_data = 12'h4a3;
			{8'd73, 8'd56}: color_data = 12'h4a3;
			{8'd73, 8'd57}: color_data = 12'h4a3;
			{8'd73, 8'd58}: color_data = 12'h4a3;
			{8'd73, 8'd59}: color_data = 12'h4a3;
			{8'd73, 8'd60}: color_data = 12'h4a3;
			{8'd73, 8'd61}: color_data = 12'h4a3;
			{8'd73, 8'd62}: color_data = 12'h4a3;
			{8'd73, 8'd63}: color_data = 12'h4a3;
			{8'd73, 8'd64}: color_data = 12'h4a3;
			{8'd73, 8'd65}: color_data = 12'h4a3;
			{8'd73, 8'd66}: color_data = 12'h4b3;
			{8'd73, 8'd67}: color_data = 12'h382;
			{8'd73, 8'd68}: color_data = 12'h000;
			{8'd73, 8'd69}: color_data = 12'h000;
			{8'd73, 8'd70}: color_data = 12'h000;
			{8'd73, 8'd71}: color_data = 12'h000;
			{8'd73, 8'd72}: color_data = 12'h000;
			{8'd73, 8'd73}: color_data = 12'h000;
			{8'd73, 8'd74}: color_data = 12'h000;
			{8'd73, 8'd100}: color_data = 12'he00;
			{8'd73, 8'd101}: color_data = 12'hf01;
			{8'd73, 8'd102}: color_data = 12'he00;
			{8'd73, 8'd103}: color_data = 12'he00;
			{8'd73, 8'd104}: color_data = 12'he00;
			{8'd73, 8'd105}: color_data = 12'he00;
			{8'd73, 8'd106}: color_data = 12'hc00;
			{8'd73, 8'd124}: color_data = 12'he01;
			{8'd73, 8'd125}: color_data = 12'he00;
			{8'd73, 8'd126}: color_data = 12'he00;
			{8'd73, 8'd127}: color_data = 12'he00;
			{8'd73, 8'd128}: color_data = 12'he00;
			{8'd73, 8'd129}: color_data = 12'he00;
			{8'd73, 8'd130}: color_data = 12'he00;
			{8'd73, 8'd131}: color_data = 12'he00;
			{8'd73, 8'd132}: color_data = 12'hf01;
			{8'd73, 8'd133}: color_data = 12'he00;
			{8'd73, 8'd138}: color_data = 12'he00;
			{8'd73, 8'd139}: color_data = 12'he00;
			{8'd73, 8'd140}: color_data = 12'he00;
			{8'd73, 8'd141}: color_data = 12'he00;
			{8'd73, 8'd142}: color_data = 12'he00;
			{8'd73, 8'd143}: color_data = 12'he01;
			{8'd73, 8'd144}: color_data = 12'he00;
			{8'd74, 8'd7}: color_data = 12'h000;
			{8'd74, 8'd8}: color_data = 12'h000;
			{8'd74, 8'd9}: color_data = 12'h000;
			{8'd74, 8'd10}: color_data = 12'ha80;
			{8'd74, 8'd11}: color_data = 12'hfd0;
			{8'd74, 8'd12}: color_data = 12'hfc0;
			{8'd74, 8'd13}: color_data = 12'hfc0;
			{8'd74, 8'd14}: color_data = 12'hfc0;
			{8'd74, 8'd15}: color_data = 12'hfc0;
			{8'd74, 8'd16}: color_data = 12'hfc0;
			{8'd74, 8'd17}: color_data = 12'hfc0;
			{8'd74, 8'd18}: color_data = 12'hfc0;
			{8'd74, 8'd19}: color_data = 12'hfc0;
			{8'd74, 8'd20}: color_data = 12'hfc0;
			{8'd74, 8'd21}: color_data = 12'hfc0;
			{8'd74, 8'd22}: color_data = 12'hfd0;
			{8'd74, 8'd23}: color_data = 12'hfd0;
			{8'd74, 8'd24}: color_data = 12'hfd0;
			{8'd74, 8'd25}: color_data = 12'hfc0;
			{8'd74, 8'd26}: color_data = 12'h540;
			{8'd74, 8'd27}: color_data = 12'h000;
			{8'd74, 8'd28}: color_data = 12'h000;
			{8'd74, 8'd29}: color_data = 12'h000;
			{8'd74, 8'd30}: color_data = 12'h000;
			{8'd74, 8'd31}: color_data = 12'h000;
			{8'd74, 8'd32}: color_data = 12'h000;
			{8'd74, 8'd33}: color_data = 12'h000;
			{8'd74, 8'd34}: color_data = 12'h000;
			{8'd74, 8'd35}: color_data = 12'h000;
			{8'd74, 8'd36}: color_data = 12'h000;
			{8'd74, 8'd37}: color_data = 12'h000;
			{8'd74, 8'd38}: color_data = 12'h000;
			{8'd74, 8'd39}: color_data = 12'h000;
			{8'd74, 8'd40}: color_data = 12'h000;
			{8'd74, 8'd41}: color_data = 12'h000;
			{8'd74, 8'd42}: color_data = 12'h130;
			{8'd74, 8'd43}: color_data = 12'h262;
			{8'd74, 8'd44}: color_data = 12'h392;
			{8'd74, 8'd45}: color_data = 12'h4b3;
			{8'd74, 8'd46}: color_data = 12'h4b3;
			{8'd74, 8'd47}: color_data = 12'h4b3;
			{8'd74, 8'd48}: color_data = 12'h4a3;
			{8'd74, 8'd49}: color_data = 12'h4a3;
			{8'd74, 8'd50}: color_data = 12'h4a3;
			{8'd74, 8'd51}: color_data = 12'h4a3;
			{8'd74, 8'd52}: color_data = 12'h4a3;
			{8'd74, 8'd53}: color_data = 12'h4a3;
			{8'd74, 8'd54}: color_data = 12'h4a3;
			{8'd74, 8'd55}: color_data = 12'h4a3;
			{8'd74, 8'd56}: color_data = 12'h4a3;
			{8'd74, 8'd57}: color_data = 12'h4a3;
			{8'd74, 8'd58}: color_data = 12'h4a3;
			{8'd74, 8'd59}: color_data = 12'h4a3;
			{8'd74, 8'd60}: color_data = 12'h4a3;
			{8'd74, 8'd61}: color_data = 12'h4a3;
			{8'd74, 8'd62}: color_data = 12'h4a3;
			{8'd74, 8'd63}: color_data = 12'h4a3;
			{8'd74, 8'd64}: color_data = 12'h4a3;
			{8'd74, 8'd65}: color_data = 12'h4a3;
			{8'd74, 8'd66}: color_data = 12'h4b3;
			{8'd74, 8'd67}: color_data = 12'h262;
			{8'd74, 8'd68}: color_data = 12'h000;
			{8'd74, 8'd69}: color_data = 12'h000;
			{8'd74, 8'd70}: color_data = 12'h000;
			{8'd74, 8'd71}: color_data = 12'h000;
			{8'd74, 8'd72}: color_data = 12'h000;
			{8'd74, 8'd73}: color_data = 12'h000;
			{8'd74, 8'd74}: color_data = 12'h000;
			{8'd74, 8'd100}: color_data = 12'he00;
			{8'd74, 8'd101}: color_data = 12'hf01;
			{8'd74, 8'd102}: color_data = 12'he00;
			{8'd74, 8'd103}: color_data = 12'he00;
			{8'd74, 8'd104}: color_data = 12'he00;
			{8'd74, 8'd105}: color_data = 12'he00;
			{8'd74, 8'd106}: color_data = 12'hc00;
			{8'd74, 8'd121}: color_data = 12'he00;
			{8'd74, 8'd122}: color_data = 12'he00;
			{8'd74, 8'd123}: color_data = 12'he00;
			{8'd74, 8'd124}: color_data = 12'he00;
			{8'd74, 8'd125}: color_data = 12'he00;
			{8'd74, 8'd126}: color_data = 12'he01;
			{8'd74, 8'd127}: color_data = 12'he00;
			{8'd74, 8'd128}: color_data = 12'he00;
			{8'd74, 8'd129}: color_data = 12'he00;
			{8'd74, 8'd130}: color_data = 12'he00;
			{8'd74, 8'd131}: color_data = 12'he00;
			{8'd74, 8'd132}: color_data = 12'hf01;
			{8'd74, 8'd133}: color_data = 12'he00;
			{8'd74, 8'd138}: color_data = 12'he00;
			{8'd74, 8'd139}: color_data = 12'he00;
			{8'd74, 8'd140}: color_data = 12'he00;
			{8'd74, 8'd141}: color_data = 12'he00;
			{8'd74, 8'd142}: color_data = 12'he00;
			{8'd74, 8'd143}: color_data = 12'he01;
			{8'd74, 8'd144}: color_data = 12'he00;
			{8'd75, 8'd4}: color_data = 12'h000;
			{8'd75, 8'd5}: color_data = 12'h000;
			{8'd75, 8'd6}: color_data = 12'h000;
			{8'd75, 8'd7}: color_data = 12'h000;
			{8'd75, 8'd8}: color_data = 12'h000;
			{8'd75, 8'd9}: color_data = 12'h000;
			{8'd75, 8'd10}: color_data = 12'h860;
			{8'd75, 8'd11}: color_data = 12'hfd0;
			{8'd75, 8'd12}: color_data = 12'hfc0;
			{8'd75, 8'd13}: color_data = 12'hfc0;
			{8'd75, 8'd14}: color_data = 12'hfc0;
			{8'd75, 8'd15}: color_data = 12'hfc0;
			{8'd75, 8'd16}: color_data = 12'hfd0;
			{8'd75, 8'd17}: color_data = 12'hfd0;
			{8'd75, 8'd18}: color_data = 12'hfd0;
			{8'd75, 8'd19}: color_data = 12'hfd0;
			{8'd75, 8'd20}: color_data = 12'hfd0;
			{8'd75, 8'd21}: color_data = 12'hfd0;
			{8'd75, 8'd22}: color_data = 12'hfc0;
			{8'd75, 8'd23}: color_data = 12'hdb0;
			{8'd75, 8'd24}: color_data = 12'hb90;
			{8'd75, 8'd25}: color_data = 12'h430;
			{8'd75, 8'd26}: color_data = 12'h000;
			{8'd75, 8'd27}: color_data = 12'h000;
			{8'd75, 8'd28}: color_data = 12'h000;
			{8'd75, 8'd29}: color_data = 12'h000;
			{8'd75, 8'd30}: color_data = 12'h000;
			{8'd75, 8'd31}: color_data = 12'h000;
			{8'd75, 8'd32}: color_data = 12'h000;
			{8'd75, 8'd33}: color_data = 12'h000;
			{8'd75, 8'd34}: color_data = 12'h000;
			{8'd75, 8'd35}: color_data = 12'h000;
			{8'd75, 8'd36}: color_data = 12'h000;
			{8'd75, 8'd37}: color_data = 12'h000;
			{8'd75, 8'd38}: color_data = 12'h000;
			{8'd75, 8'd39}: color_data = 12'h000;
			{8'd75, 8'd40}: color_data = 12'h000;
			{8'd75, 8'd41}: color_data = 12'h000;
			{8'd75, 8'd42}: color_data = 12'h000;
			{8'd75, 8'd43}: color_data = 12'h000;
			{8'd75, 8'd44}: color_data = 12'h000;
			{8'd75, 8'd45}: color_data = 12'h131;
			{8'd75, 8'd46}: color_data = 12'h272;
			{8'd75, 8'd47}: color_data = 12'h3a3;
			{8'd75, 8'd48}: color_data = 12'h4b3;
			{8'd75, 8'd49}: color_data = 12'h4b3;
			{8'd75, 8'd50}: color_data = 12'h4b3;
			{8'd75, 8'd51}: color_data = 12'h4a3;
			{8'd75, 8'd52}: color_data = 12'h4a3;
			{8'd75, 8'd53}: color_data = 12'h4a3;
			{8'd75, 8'd54}: color_data = 12'h4a3;
			{8'd75, 8'd55}: color_data = 12'h4a3;
			{8'd75, 8'd56}: color_data = 12'h4a3;
			{8'd75, 8'd57}: color_data = 12'h4a3;
			{8'd75, 8'd58}: color_data = 12'h4a3;
			{8'd75, 8'd59}: color_data = 12'h4a3;
			{8'd75, 8'd60}: color_data = 12'h4a3;
			{8'd75, 8'd61}: color_data = 12'h4a3;
			{8'd75, 8'd62}: color_data = 12'h4a3;
			{8'd75, 8'd63}: color_data = 12'h4a3;
			{8'd75, 8'd64}: color_data = 12'h4a3;
			{8'd75, 8'd65}: color_data = 12'h4a3;
			{8'd75, 8'd66}: color_data = 12'h4b3;
			{8'd75, 8'd67}: color_data = 12'h141;
			{8'd75, 8'd68}: color_data = 12'h000;
			{8'd75, 8'd69}: color_data = 12'h000;
			{8'd75, 8'd70}: color_data = 12'h000;
			{8'd75, 8'd71}: color_data = 12'h000;
			{8'd75, 8'd72}: color_data = 12'h000;
			{8'd75, 8'd73}: color_data = 12'h000;
			{8'd75, 8'd74}: color_data = 12'h000;
			{8'd75, 8'd100}: color_data = 12'he00;
			{8'd75, 8'd101}: color_data = 12'hf01;
			{8'd75, 8'd102}: color_data = 12'he00;
			{8'd75, 8'd103}: color_data = 12'he00;
			{8'd75, 8'd104}: color_data = 12'he00;
			{8'd75, 8'd105}: color_data = 12'he00;
			{8'd75, 8'd106}: color_data = 12'hc00;
			{8'd75, 8'd117}: color_data = 12'hf00;
			{8'd75, 8'd118}: color_data = 12'he00;
			{8'd75, 8'd119}: color_data = 12'he00;
			{8'd75, 8'd120}: color_data = 12'he00;
			{8'd75, 8'd121}: color_data = 12'he00;
			{8'd75, 8'd122}: color_data = 12'he01;
			{8'd75, 8'd123}: color_data = 12'he01;
			{8'd75, 8'd124}: color_data = 12'he00;
			{8'd75, 8'd125}: color_data = 12'he00;
			{8'd75, 8'd126}: color_data = 12'he00;
			{8'd75, 8'd127}: color_data = 12'he00;
			{8'd75, 8'd128}: color_data = 12'he00;
			{8'd75, 8'd129}: color_data = 12'he00;
			{8'd75, 8'd130}: color_data = 12'he00;
			{8'd75, 8'd131}: color_data = 12'he01;
			{8'd75, 8'd132}: color_data = 12'he00;
			{8'd75, 8'd133}: color_data = 12'he00;
			{8'd75, 8'd138}: color_data = 12'he00;
			{8'd75, 8'd139}: color_data = 12'he00;
			{8'd75, 8'd140}: color_data = 12'he00;
			{8'd75, 8'd141}: color_data = 12'he00;
			{8'd75, 8'd142}: color_data = 12'he00;
			{8'd75, 8'd143}: color_data = 12'he01;
			{8'd75, 8'd144}: color_data = 12'he00;
			{8'd76, 8'd4}: color_data = 12'h000;
			{8'd76, 8'd5}: color_data = 12'h000;
			{8'd76, 8'd6}: color_data = 12'h000;
			{8'd76, 8'd7}: color_data = 12'h000;
			{8'd76, 8'd8}: color_data = 12'h000;
			{8'd76, 8'd9}: color_data = 12'h000;
			{8'd76, 8'd10}: color_data = 12'h650;
			{8'd76, 8'd11}: color_data = 12'hfd0;
			{8'd76, 8'd12}: color_data = 12'hfd0;
			{8'd76, 8'd13}: color_data = 12'hfd0;
			{8'd76, 8'd14}: color_data = 12'hfd0;
			{8'd76, 8'd15}: color_data = 12'hfd0;
			{8'd76, 8'd16}: color_data = 12'hfc0;
			{8'd76, 8'd17}: color_data = 12'hdb0;
			{8'd76, 8'd18}: color_data = 12'hb90;
			{8'd76, 8'd19}: color_data = 12'h970;
			{8'd76, 8'd20}: color_data = 12'h650;
			{8'd76, 8'd21}: color_data = 12'h430;
			{8'd76, 8'd22}: color_data = 12'h210;
			{8'd76, 8'd23}: color_data = 12'h000;
			{8'd76, 8'd24}: color_data = 12'h000;
			{8'd76, 8'd25}: color_data = 12'h000;
			{8'd76, 8'd26}: color_data = 12'h000;
			{8'd76, 8'd27}: color_data = 12'h000;
			{8'd76, 8'd28}: color_data = 12'h000;
			{8'd76, 8'd29}: color_data = 12'h000;
			{8'd76, 8'd30}: color_data = 12'h000;
			{8'd76, 8'd31}: color_data = 12'h000;
			{8'd76, 8'd32}: color_data = 12'h000;
			{8'd76, 8'd33}: color_data = 12'h000;
			{8'd76, 8'd34}: color_data = 12'h000;
			{8'd76, 8'd35}: color_data = 12'h000;
			{8'd76, 8'd36}: color_data = 12'h000;
			{8'd76, 8'd37}: color_data = 12'h000;
			{8'd76, 8'd38}: color_data = 12'h000;
			{8'd76, 8'd39}: color_data = 12'h000;
			{8'd76, 8'd40}: color_data = 12'h000;
			{8'd76, 8'd41}: color_data = 12'h000;
			{8'd76, 8'd42}: color_data = 12'h000;
			{8'd76, 8'd43}: color_data = 12'h000;
			{8'd76, 8'd44}: color_data = 12'h000;
			{8'd76, 8'd45}: color_data = 12'h000;
			{8'd76, 8'd46}: color_data = 12'h000;
			{8'd76, 8'd47}: color_data = 12'h010;
			{8'd76, 8'd48}: color_data = 12'h131;
			{8'd76, 8'd49}: color_data = 12'h272;
			{8'd76, 8'd50}: color_data = 12'h4a3;
			{8'd76, 8'd51}: color_data = 12'h4b3;
			{8'd76, 8'd52}: color_data = 12'h4b3;
			{8'd76, 8'd53}: color_data = 12'h4b3;
			{8'd76, 8'd54}: color_data = 12'h4a3;
			{8'd76, 8'd55}: color_data = 12'h4a3;
			{8'd76, 8'd56}: color_data = 12'h4a3;
			{8'd76, 8'd57}: color_data = 12'h4a3;
			{8'd76, 8'd58}: color_data = 12'h4a3;
			{8'd76, 8'd59}: color_data = 12'h4a3;
			{8'd76, 8'd60}: color_data = 12'h4a3;
			{8'd76, 8'd61}: color_data = 12'h4a3;
			{8'd76, 8'd62}: color_data = 12'h4a3;
			{8'd76, 8'd63}: color_data = 12'h4a3;
			{8'd76, 8'd64}: color_data = 12'h4a3;
			{8'd76, 8'd65}: color_data = 12'h4b3;
			{8'd76, 8'd66}: color_data = 12'h4b3;
			{8'd76, 8'd67}: color_data = 12'h120;
			{8'd76, 8'd68}: color_data = 12'h000;
			{8'd76, 8'd69}: color_data = 12'h000;
			{8'd76, 8'd70}: color_data = 12'h000;
			{8'd76, 8'd71}: color_data = 12'h000;
			{8'd76, 8'd72}: color_data = 12'h000;
			{8'd76, 8'd73}: color_data = 12'h000;
			{8'd76, 8'd74}: color_data = 12'h000;
			{8'd76, 8'd100}: color_data = 12'he00;
			{8'd76, 8'd101}: color_data = 12'hf01;
			{8'd76, 8'd102}: color_data = 12'he00;
			{8'd76, 8'd103}: color_data = 12'he00;
			{8'd76, 8'd104}: color_data = 12'he00;
			{8'd76, 8'd105}: color_data = 12'he00;
			{8'd76, 8'd106}: color_data = 12'hc00;
			{8'd76, 8'd117}: color_data = 12'he00;
			{8'd76, 8'd118}: color_data = 12'he00;
			{8'd76, 8'd119}: color_data = 12'he01;
			{8'd76, 8'd120}: color_data = 12'he01;
			{8'd76, 8'd121}: color_data = 12'he00;
			{8'd76, 8'd122}: color_data = 12'he00;
			{8'd76, 8'd123}: color_data = 12'he00;
			{8'd76, 8'd124}: color_data = 12'he00;
			{8'd76, 8'd125}: color_data = 12'he00;
			{8'd76, 8'd126}: color_data = 12'he00;
			{8'd76, 8'd127}: color_data = 12'he00;
			{8'd76, 8'd128}: color_data = 12'he00;
			{8'd76, 8'd129}: color_data = 12'he00;
			{8'd76, 8'd130}: color_data = 12'he00;
			{8'd76, 8'd131}: color_data = 12'he00;
			{8'd76, 8'd132}: color_data = 12'he00;
			{8'd76, 8'd138}: color_data = 12'he00;
			{8'd76, 8'd139}: color_data = 12'he00;
			{8'd76, 8'd140}: color_data = 12'he00;
			{8'd76, 8'd141}: color_data = 12'he00;
			{8'd76, 8'd142}: color_data = 12'he00;
			{8'd76, 8'd143}: color_data = 12'he01;
			{8'd76, 8'd144}: color_data = 12'he00;
			{8'd77, 8'd4}: color_data = 12'h000;
			{8'd77, 8'd5}: color_data = 12'h000;
			{8'd77, 8'd6}: color_data = 12'h000;
			{8'd77, 8'd7}: color_data = 12'h000;
			{8'd77, 8'd8}: color_data = 12'h000;
			{8'd77, 8'd9}: color_data = 12'h000;
			{8'd77, 8'd10}: color_data = 12'h330;
			{8'd77, 8'd11}: color_data = 12'hdb0;
			{8'd77, 8'd12}: color_data = 12'hb90;
			{8'd77, 8'd13}: color_data = 12'h970;
			{8'd77, 8'd14}: color_data = 12'h650;
			{8'd77, 8'd15}: color_data = 12'h430;
			{8'd77, 8'd16}: color_data = 12'h210;
			{8'd77, 8'd17}: color_data = 12'h000;
			{8'd77, 8'd18}: color_data = 12'h000;
			{8'd77, 8'd19}: color_data = 12'h000;
			{8'd77, 8'd20}: color_data = 12'h000;
			{8'd77, 8'd21}: color_data = 12'h000;
			{8'd77, 8'd22}: color_data = 12'h000;
			{8'd77, 8'd23}: color_data = 12'h000;
			{8'd77, 8'd24}: color_data = 12'h000;
			{8'd77, 8'd25}: color_data = 12'h000;
			{8'd77, 8'd26}: color_data = 12'h000;
			{8'd77, 8'd27}: color_data = 12'h000;
			{8'd77, 8'd28}: color_data = 12'h000;
			{8'd77, 8'd29}: color_data = 12'h000;
			{8'd77, 8'd30}: color_data = 12'h000;
			{8'd77, 8'd31}: color_data = 12'h000;
			{8'd77, 8'd32}: color_data = 12'h000;
			{8'd77, 8'd33}: color_data = 12'h000;
			{8'd77, 8'd34}: color_data = 12'h000;
			{8'd77, 8'd35}: color_data = 12'h000;
			{8'd77, 8'd36}: color_data = 12'h000;
			{8'd77, 8'd37}: color_data = 12'h000;
			{8'd77, 8'd38}: color_data = 12'h000;
			{8'd77, 8'd39}: color_data = 12'h000;
			{8'd77, 8'd40}: color_data = 12'h000;
			{8'd77, 8'd41}: color_data = 12'h000;
			{8'd77, 8'd42}: color_data = 12'h000;
			{8'd77, 8'd43}: color_data = 12'h000;
			{8'd77, 8'd44}: color_data = 12'h000;
			{8'd77, 8'd45}: color_data = 12'h000;
			{8'd77, 8'd46}: color_data = 12'h000;
			{8'd77, 8'd47}: color_data = 12'h000;
			{8'd77, 8'd48}: color_data = 12'h000;
			{8'd77, 8'd49}: color_data = 12'h000;
			{8'd77, 8'd50}: color_data = 12'h010;
			{8'd77, 8'd51}: color_data = 12'h141;
			{8'd77, 8'd52}: color_data = 12'h382;
			{8'd77, 8'd53}: color_data = 12'h4a3;
			{8'd77, 8'd54}: color_data = 12'h4b3;
			{8'd77, 8'd55}: color_data = 12'h4b3;
			{8'd77, 8'd56}: color_data = 12'h4b3;
			{8'd77, 8'd57}: color_data = 12'h4a3;
			{8'd77, 8'd58}: color_data = 12'h4a3;
			{8'd77, 8'd59}: color_data = 12'h4a3;
			{8'd77, 8'd60}: color_data = 12'h4a3;
			{8'd77, 8'd61}: color_data = 12'h4a3;
			{8'd77, 8'd62}: color_data = 12'h4a3;
			{8'd77, 8'd63}: color_data = 12'h4a3;
			{8'd77, 8'd64}: color_data = 12'h4a3;
			{8'd77, 8'd65}: color_data = 12'h4b3;
			{8'd77, 8'd66}: color_data = 12'h4a3;
			{8'd77, 8'd67}: color_data = 12'h010;
			{8'd77, 8'd68}: color_data = 12'h000;
			{8'd77, 8'd69}: color_data = 12'h000;
			{8'd77, 8'd70}: color_data = 12'h000;
			{8'd77, 8'd71}: color_data = 12'h000;
			{8'd77, 8'd72}: color_data = 12'h000;
			{8'd77, 8'd73}: color_data = 12'h000;
			{8'd77, 8'd74}: color_data = 12'h000;
			{8'd77, 8'd100}: color_data = 12'he00;
			{8'd77, 8'd101}: color_data = 12'hf01;
			{8'd77, 8'd102}: color_data = 12'he00;
			{8'd77, 8'd103}: color_data = 12'he00;
			{8'd77, 8'd104}: color_data = 12'he00;
			{8'd77, 8'd105}: color_data = 12'he00;
			{8'd77, 8'd106}: color_data = 12'hc00;
			{8'd77, 8'd117}: color_data = 12'he00;
			{8'd77, 8'd118}: color_data = 12'he00;
			{8'd77, 8'd119}: color_data = 12'he00;
			{8'd77, 8'd120}: color_data = 12'he00;
			{8'd77, 8'd121}: color_data = 12'he00;
			{8'd77, 8'd122}: color_data = 12'he00;
			{8'd77, 8'd123}: color_data = 12'he00;
			{8'd77, 8'd124}: color_data = 12'he00;
			{8'd77, 8'd125}: color_data = 12'he00;
			{8'd77, 8'd126}: color_data = 12'hf01;
			{8'd77, 8'd127}: color_data = 12'he00;
			{8'd77, 8'd128}: color_data = 12'he00;
			{8'd77, 8'd129}: color_data = 12'he00;
			{8'd77, 8'd130}: color_data = 12'hf00;
			{8'd77, 8'd138}: color_data = 12'he00;
			{8'd77, 8'd139}: color_data = 12'he00;
			{8'd77, 8'd140}: color_data = 12'he00;
			{8'd77, 8'd141}: color_data = 12'he00;
			{8'd77, 8'd142}: color_data = 12'he00;
			{8'd77, 8'd143}: color_data = 12'he01;
			{8'd77, 8'd144}: color_data = 12'he00;
			{8'd78, 8'd4}: color_data = 12'h000;
			{8'd78, 8'd5}: color_data = 12'h000;
			{8'd78, 8'd6}: color_data = 12'h300;
			{8'd78, 8'd7}: color_data = 12'h810;
			{8'd78, 8'd8}: color_data = 12'h400;
			{8'd78, 8'd9}: color_data = 12'h000;
			{8'd78, 8'd10}: color_data = 12'h000;
			{8'd78, 8'd11}: color_data = 12'h000;
			{8'd78, 8'd12}: color_data = 12'h000;
			{8'd78, 8'd13}: color_data = 12'h000;
			{8'd78, 8'd14}: color_data = 12'h000;
			{8'd78, 8'd15}: color_data = 12'h000;
			{8'd78, 8'd16}: color_data = 12'h000;
			{8'd78, 8'd17}: color_data = 12'h000;
			{8'd78, 8'd18}: color_data = 12'h000;
			{8'd78, 8'd19}: color_data = 12'h000;
			{8'd78, 8'd20}: color_data = 12'h000;
			{8'd78, 8'd21}: color_data = 12'h000;
			{8'd78, 8'd22}: color_data = 12'h000;
			{8'd78, 8'd23}: color_data = 12'h000;
			{8'd78, 8'd24}: color_data = 12'h000;
			{8'd78, 8'd25}: color_data = 12'h000;
			{8'd78, 8'd26}: color_data = 12'h000;
			{8'd78, 8'd27}: color_data = 12'h000;
			{8'd78, 8'd28}: color_data = 12'h000;
			{8'd78, 8'd29}: color_data = 12'h000;
			{8'd78, 8'd30}: color_data = 12'h000;
			{8'd78, 8'd31}: color_data = 12'h000;
			{8'd78, 8'd32}: color_data = 12'h000;
			{8'd78, 8'd33}: color_data = 12'h000;
			{8'd78, 8'd34}: color_data = 12'h000;
			{8'd78, 8'd35}: color_data = 12'h000;
			{8'd78, 8'd36}: color_data = 12'h000;
			{8'd78, 8'd37}: color_data = 12'h000;
			{8'd78, 8'd38}: color_data = 12'h000;
			{8'd78, 8'd39}: color_data = 12'h000;
			{8'd78, 8'd40}: color_data = 12'h000;
			{8'd78, 8'd41}: color_data = 12'h000;
			{8'd78, 8'd42}: color_data = 12'h000;
			{8'd78, 8'd43}: color_data = 12'h000;
			{8'd78, 8'd44}: color_data = 12'h000;
			{8'd78, 8'd45}: color_data = 12'h000;
			{8'd78, 8'd46}: color_data = 12'h000;
			{8'd78, 8'd47}: color_data = 12'h000;
			{8'd78, 8'd48}: color_data = 12'h000;
			{8'd78, 8'd49}: color_data = 12'h000;
			{8'd78, 8'd50}: color_data = 12'h000;
			{8'd78, 8'd51}: color_data = 12'h000;
			{8'd78, 8'd52}: color_data = 12'h000;
			{8'd78, 8'd53}: color_data = 12'h010;
			{8'd78, 8'd54}: color_data = 12'h141;
			{8'd78, 8'd55}: color_data = 12'h382;
			{8'd78, 8'd56}: color_data = 12'h4a3;
			{8'd78, 8'd57}: color_data = 12'h4b3;
			{8'd78, 8'd58}: color_data = 12'h4b3;
			{8'd78, 8'd59}: color_data = 12'h4b3;
			{8'd78, 8'd60}: color_data = 12'h4a3;
			{8'd78, 8'd61}: color_data = 12'h4a3;
			{8'd78, 8'd62}: color_data = 12'h4a3;
			{8'd78, 8'd63}: color_data = 12'h4a3;
			{8'd78, 8'd64}: color_data = 12'h4a3;
			{8'd78, 8'd65}: color_data = 12'h4b3;
			{8'd78, 8'd66}: color_data = 12'h392;
			{8'd78, 8'd67}: color_data = 12'h000;
			{8'd78, 8'd68}: color_data = 12'h000;
			{8'd78, 8'd69}: color_data = 12'h000;
			{8'd78, 8'd70}: color_data = 12'h000;
			{8'd78, 8'd71}: color_data = 12'h000;
			{8'd78, 8'd72}: color_data = 12'h000;
			{8'd78, 8'd73}: color_data = 12'h000;
			{8'd78, 8'd100}: color_data = 12'he00;
			{8'd78, 8'd101}: color_data = 12'hf01;
			{8'd78, 8'd102}: color_data = 12'he00;
			{8'd78, 8'd103}: color_data = 12'he00;
			{8'd78, 8'd104}: color_data = 12'he00;
			{8'd78, 8'd105}: color_data = 12'he00;
			{8'd78, 8'd106}: color_data = 12'hc00;
			{8'd78, 8'd117}: color_data = 12'he00;
			{8'd78, 8'd118}: color_data = 12'he00;
			{8'd78, 8'd119}: color_data = 12'he00;
			{8'd78, 8'd120}: color_data = 12'he00;
			{8'd78, 8'd121}: color_data = 12'he00;
			{8'd78, 8'd122}: color_data = 12'he00;
			{8'd78, 8'd123}: color_data = 12'he00;
			{8'd78, 8'd124}: color_data = 12'he01;
			{8'd78, 8'd125}: color_data = 12'he00;
			{8'd78, 8'd126}: color_data = 12'he01;
			{8'd78, 8'd127}: color_data = 12'he00;
			{8'd78, 8'd138}: color_data = 12'he00;
			{8'd78, 8'd139}: color_data = 12'he00;
			{8'd78, 8'd140}: color_data = 12'he00;
			{8'd78, 8'd141}: color_data = 12'he00;
			{8'd78, 8'd142}: color_data = 12'he00;
			{8'd78, 8'd143}: color_data = 12'he01;
			{8'd78, 8'd144}: color_data = 12'he00;
			{8'd79, 8'd3}: color_data = 12'h000;
			{8'd79, 8'd4}: color_data = 12'h000;
			{8'd79, 8'd5}: color_data = 12'h000;
			{8'd79, 8'd6}: color_data = 12'h710;
			{8'd79, 8'd7}: color_data = 12'hf21;
			{8'd79, 8'd8}: color_data = 12'ha10;
			{8'd79, 8'd9}: color_data = 12'h000;
			{8'd79, 8'd10}: color_data = 12'h000;
			{8'd79, 8'd11}: color_data = 12'h000;
			{8'd79, 8'd12}: color_data = 12'h000;
			{8'd79, 8'd13}: color_data = 12'h200;
			{8'd79, 8'd14}: color_data = 12'h400;
			{8'd79, 8'd15}: color_data = 12'h610;
			{8'd79, 8'd16}: color_data = 12'h710;
			{8'd79, 8'd17}: color_data = 12'h500;
			{8'd79, 8'd18}: color_data = 12'h300;
			{8'd79, 8'd19}: color_data = 12'h200;
			{8'd79, 8'd20}: color_data = 12'h100;
			{8'd79, 8'd21}: color_data = 12'h000;
			{8'd79, 8'd22}: color_data = 12'h000;
			{8'd79, 8'd23}: color_data = 12'h000;
			{8'd79, 8'd24}: color_data = 12'h000;
			{8'd79, 8'd25}: color_data = 12'h000;
			{8'd79, 8'd26}: color_data = 12'h000;
			{8'd79, 8'd27}: color_data = 12'h000;
			{8'd79, 8'd28}: color_data = 12'h000;
			{8'd79, 8'd29}: color_data = 12'h000;
			{8'd79, 8'd30}: color_data = 12'h000;
			{8'd79, 8'd31}: color_data = 12'h000;
			{8'd79, 8'd32}: color_data = 12'h000;
			{8'd79, 8'd33}: color_data = 12'h000;
			{8'd79, 8'd34}: color_data = 12'h000;
			{8'd79, 8'd35}: color_data = 12'h110;
			{8'd79, 8'd36}: color_data = 12'h650;
			{8'd79, 8'd37}: color_data = 12'h440;
			{8'd79, 8'd38}: color_data = 12'h320;
			{8'd79, 8'd39}: color_data = 12'h110;
			{8'd79, 8'd40}: color_data = 12'h000;
			{8'd79, 8'd41}: color_data = 12'h000;
			{8'd79, 8'd42}: color_data = 12'h000;
			{8'd79, 8'd43}: color_data = 12'h000;
			{8'd79, 8'd44}: color_data = 12'h000;
			{8'd79, 8'd45}: color_data = 12'h000;
			{8'd79, 8'd46}: color_data = 12'h000;
			{8'd79, 8'd47}: color_data = 12'h000;
			{8'd79, 8'd48}: color_data = 12'h000;
			{8'd79, 8'd49}: color_data = 12'h000;
			{8'd79, 8'd50}: color_data = 12'h000;
			{8'd79, 8'd51}: color_data = 12'h000;
			{8'd79, 8'd52}: color_data = 12'h000;
			{8'd79, 8'd53}: color_data = 12'h000;
			{8'd79, 8'd54}: color_data = 12'h000;
			{8'd79, 8'd55}: color_data = 12'h000;
			{8'd79, 8'd56}: color_data = 12'h010;
			{8'd79, 8'd57}: color_data = 12'h251;
			{8'd79, 8'd58}: color_data = 12'h382;
			{8'd79, 8'd59}: color_data = 12'h4a3;
			{8'd79, 8'd60}: color_data = 12'h4b3;
			{8'd79, 8'd61}: color_data = 12'h4b3;
			{8'd79, 8'd62}: color_data = 12'h4b3;
			{8'd79, 8'd63}: color_data = 12'h4a3;
			{8'd79, 8'd64}: color_data = 12'h4a3;
			{8'd79, 8'd65}: color_data = 12'h4b3;
			{8'd79, 8'd66}: color_data = 12'h272;
			{8'd79, 8'd67}: color_data = 12'h000;
			{8'd79, 8'd68}: color_data = 12'h000;
			{8'd79, 8'd69}: color_data = 12'h000;
			{8'd79, 8'd70}: color_data = 12'h000;
			{8'd79, 8'd71}: color_data = 12'h000;
			{8'd79, 8'd72}: color_data = 12'h000;
			{8'd79, 8'd73}: color_data = 12'h000;
			{8'd79, 8'd100}: color_data = 12'he00;
			{8'd79, 8'd101}: color_data = 12'hf01;
			{8'd79, 8'd102}: color_data = 12'he00;
			{8'd79, 8'd103}: color_data = 12'he00;
			{8'd79, 8'd104}: color_data = 12'he00;
			{8'd79, 8'd105}: color_data = 12'he00;
			{8'd79, 8'd106}: color_data = 12'hc00;
			{8'd79, 8'd117}: color_data = 12'he00;
			{8'd79, 8'd118}: color_data = 12'he00;
			{8'd79, 8'd119}: color_data = 12'he00;
			{8'd79, 8'd120}: color_data = 12'he00;
			{8'd79, 8'd121}: color_data = 12'he01;
			{8'd79, 8'd122}: color_data = 12'he00;
			{8'd79, 8'd123}: color_data = 12'he00;
			{8'd79, 8'd124}: color_data = 12'he00;
			{8'd79, 8'd125}: color_data = 12'he00;
			{8'd79, 8'd138}: color_data = 12'he00;
			{8'd79, 8'd139}: color_data = 12'he00;
			{8'd79, 8'd140}: color_data = 12'he00;
			{8'd79, 8'd141}: color_data = 12'he00;
			{8'd79, 8'd142}: color_data = 12'he00;
			{8'd79, 8'd143}: color_data = 12'he01;
			{8'd79, 8'd144}: color_data = 12'he00;
			{8'd80, 8'd3}: color_data = 12'h000;
			{8'd80, 8'd4}: color_data = 12'h000;
			{8'd80, 8'd5}: color_data = 12'h000;
			{8'd80, 8'd6}: color_data = 12'ha10;
			{8'd80, 8'd7}: color_data = 12'hf21;
			{8'd80, 8'd8}: color_data = 12'hd20;
			{8'd80, 8'd9}: color_data = 12'h710;
			{8'd80, 8'd10}: color_data = 12'h810;
			{8'd80, 8'd11}: color_data = 12'hb10;
			{8'd80, 8'd12}: color_data = 12'hc10;
			{8'd80, 8'd13}: color_data = 12'he21;
			{8'd80, 8'd14}: color_data = 12'he21;
			{8'd80, 8'd15}: color_data = 12'he21;
			{8'd80, 8'd16}: color_data = 12'he21;
			{8'd80, 8'd17}: color_data = 12'he21;
			{8'd80, 8'd18}: color_data = 12'he21;
			{8'd80, 8'd19}: color_data = 12'he21;
			{8'd80, 8'd20}: color_data = 12'hd20;
			{8'd80, 8'd21}: color_data = 12'hc10;
			{8'd80, 8'd22}: color_data = 12'ha10;
			{8'd80, 8'd23}: color_data = 12'h910;
			{8'd80, 8'd24}: color_data = 12'h710;
			{8'd80, 8'd25}: color_data = 12'h500;
			{8'd80, 8'd26}: color_data = 12'h400;
			{8'd80, 8'd27}: color_data = 12'h200;
			{8'd80, 8'd28}: color_data = 12'h100;
			{8'd80, 8'd29}: color_data = 12'h000;
			{8'd80, 8'd30}: color_data = 12'h000;
			{8'd80, 8'd31}: color_data = 12'h000;
			{8'd80, 8'd32}: color_data = 12'h000;
			{8'd80, 8'd33}: color_data = 12'h000;
			{8'd80, 8'd34}: color_data = 12'h000;
			{8'd80, 8'd35}: color_data = 12'h540;
			{8'd80, 8'd36}: color_data = 12'hfd0;
			{8'd80, 8'd37}: color_data = 12'hfd0;
			{8'd80, 8'd38}: color_data = 12'hfc0;
			{8'd80, 8'd39}: color_data = 12'hec0;
			{8'd80, 8'd40}: color_data = 12'hdb0;
			{8'd80, 8'd41}: color_data = 12'hca0;
			{8'd80, 8'd42}: color_data = 12'hb90;
			{8'd80, 8'd43}: color_data = 12'h970;
			{8'd80, 8'd44}: color_data = 12'h760;
			{8'd80, 8'd45}: color_data = 12'h540;
			{8'd80, 8'd46}: color_data = 12'h430;
			{8'd80, 8'd47}: color_data = 12'h220;
			{8'd80, 8'd48}: color_data = 12'h110;
			{8'd80, 8'd49}: color_data = 12'h000;
			{8'd80, 8'd50}: color_data = 12'h000;
			{8'd80, 8'd51}: color_data = 12'h000;
			{8'd80, 8'd52}: color_data = 12'h000;
			{8'd80, 8'd53}: color_data = 12'h000;
			{8'd80, 8'd54}: color_data = 12'h000;
			{8'd80, 8'd55}: color_data = 12'h000;
			{8'd80, 8'd56}: color_data = 12'h000;
			{8'd80, 8'd57}: color_data = 12'h000;
			{8'd80, 8'd58}: color_data = 12'h000;
			{8'd80, 8'd59}: color_data = 12'h020;
			{8'd80, 8'd60}: color_data = 12'h251;
			{8'd80, 8'd61}: color_data = 12'h392;
			{8'd80, 8'd62}: color_data = 12'h4b3;
			{8'd80, 8'd63}: color_data = 12'h4b3;
			{8'd80, 8'd64}: color_data = 12'h4b3;
			{8'd80, 8'd65}: color_data = 12'h4b3;
			{8'd80, 8'd66}: color_data = 12'h251;
			{8'd80, 8'd67}: color_data = 12'h000;
			{8'd80, 8'd68}: color_data = 12'h000;
			{8'd80, 8'd69}: color_data = 12'h000;
			{8'd80, 8'd70}: color_data = 12'h000;
			{8'd80, 8'd71}: color_data = 12'h000;
			{8'd80, 8'd72}: color_data = 12'h000;
			{8'd80, 8'd73}: color_data = 12'h000;
			{8'd80, 8'd74}: color_data = 12'h000;
			{8'd80, 8'd75}: color_data = 12'h000;
			{8'd80, 8'd100}: color_data = 12'he00;
			{8'd80, 8'd101}: color_data = 12'hf01;
			{8'd80, 8'd102}: color_data = 12'he00;
			{8'd80, 8'd103}: color_data = 12'he00;
			{8'd80, 8'd104}: color_data = 12'he00;
			{8'd80, 8'd105}: color_data = 12'he00;
			{8'd80, 8'd106}: color_data = 12'hc00;
			{8'd80, 8'd117}: color_data = 12'he00;
			{8'd80, 8'd118}: color_data = 12'he00;
			{8'd80, 8'd119}: color_data = 12'hf01;
			{8'd80, 8'd120}: color_data = 12'he00;
			{8'd80, 8'd121}: color_data = 12'he00;
			{8'd80, 8'd122}: color_data = 12'he00;
			{8'd80, 8'd123}: color_data = 12'hd00;
			{8'd80, 8'd138}: color_data = 12'he00;
			{8'd80, 8'd139}: color_data = 12'he00;
			{8'd80, 8'd140}: color_data = 12'he00;
			{8'd80, 8'd141}: color_data = 12'he00;
			{8'd80, 8'd142}: color_data = 12'he00;
			{8'd80, 8'd143}: color_data = 12'he01;
			{8'd80, 8'd144}: color_data = 12'he00;
			{8'd81, 8'd3}: color_data = 12'h000;
			{8'd81, 8'd4}: color_data = 12'h000;
			{8'd81, 8'd5}: color_data = 12'h000;
			{8'd81, 8'd6}: color_data = 12'hc10;
			{8'd81, 8'd7}: color_data = 12'he21;
			{8'd81, 8'd8}: color_data = 12'he21;
			{8'd81, 8'd9}: color_data = 12'he21;
			{8'd81, 8'd10}: color_data = 12'he21;
			{8'd81, 8'd11}: color_data = 12'he21;
			{8'd81, 8'd12}: color_data = 12'he21;
			{8'd81, 8'd13}: color_data = 12'he21;
			{8'd81, 8'd14}: color_data = 12'he21;
			{8'd81, 8'd15}: color_data = 12'he21;
			{8'd81, 8'd16}: color_data = 12'he21;
			{8'd81, 8'd17}: color_data = 12'he21;
			{8'd81, 8'd18}: color_data = 12'he21;
			{8'd81, 8'd19}: color_data = 12'he21;
			{8'd81, 8'd20}: color_data = 12'he21;
			{8'd81, 8'd21}: color_data = 12'he21;
			{8'd81, 8'd22}: color_data = 12'he21;
			{8'd81, 8'd23}: color_data = 12'he21;
			{8'd81, 8'd24}: color_data = 12'hf21;
			{8'd81, 8'd25}: color_data = 12'he21;
			{8'd81, 8'd26}: color_data = 12'he21;
			{8'd81, 8'd27}: color_data = 12'he21;
			{8'd81, 8'd28}: color_data = 12'hd20;
			{8'd81, 8'd29}: color_data = 12'hc10;
			{8'd81, 8'd30}: color_data = 12'h710;
			{8'd81, 8'd31}: color_data = 12'h000;
			{8'd81, 8'd32}: color_data = 12'h000;
			{8'd81, 8'd33}: color_data = 12'h000;
			{8'd81, 8'd34}: color_data = 12'h000;
			{8'd81, 8'd35}: color_data = 12'h760;
			{8'd81, 8'd36}: color_data = 12'hfd0;
			{8'd81, 8'd37}: color_data = 12'hfc0;
			{8'd81, 8'd38}: color_data = 12'hfd0;
			{8'd81, 8'd39}: color_data = 12'hfd0;
			{8'd81, 8'd40}: color_data = 12'hfd0;
			{8'd81, 8'd41}: color_data = 12'hfd0;
			{8'd81, 8'd42}: color_data = 12'hfd0;
			{8'd81, 8'd43}: color_data = 12'hfd0;
			{8'd81, 8'd44}: color_data = 12'hfd0;
			{8'd81, 8'd45}: color_data = 12'hfd0;
			{8'd81, 8'd46}: color_data = 12'hfd0;
			{8'd81, 8'd47}: color_data = 12'hfc0;
			{8'd81, 8'd48}: color_data = 12'hec0;
			{8'd81, 8'd49}: color_data = 12'hdb0;
			{8'd81, 8'd50}: color_data = 12'hc90;
			{8'd81, 8'd51}: color_data = 12'ha80;
			{8'd81, 8'd52}: color_data = 12'h870;
			{8'd81, 8'd53}: color_data = 12'h650;
			{8'd81, 8'd54}: color_data = 12'h540;
			{8'd81, 8'd55}: color_data = 12'h330;
			{8'd81, 8'd56}: color_data = 12'h110;
			{8'd81, 8'd57}: color_data = 12'h000;
			{8'd81, 8'd58}: color_data = 12'h000;
			{8'd81, 8'd59}: color_data = 12'h000;
			{8'd81, 8'd60}: color_data = 12'h000;
			{8'd81, 8'd61}: color_data = 12'h000;
			{8'd81, 8'd62}: color_data = 12'h120;
			{8'd81, 8'd63}: color_data = 12'h261;
			{8'd81, 8'd64}: color_data = 12'h392;
			{8'd81, 8'd65}: color_data = 12'h4b3;
			{8'd81, 8'd66}: color_data = 12'h131;
			{8'd81, 8'd67}: color_data = 12'h000;
			{8'd81, 8'd68}: color_data = 12'h000;
			{8'd81, 8'd69}: color_data = 12'h000;
			{8'd81, 8'd70}: color_data = 12'h000;
			{8'd81, 8'd71}: color_data = 12'h000;
			{8'd81, 8'd72}: color_data = 12'h000;
			{8'd81, 8'd73}: color_data = 12'h000;
			{8'd81, 8'd74}: color_data = 12'h000;
			{8'd81, 8'd75}: color_data = 12'h000;
			{8'd81, 8'd100}: color_data = 12'he00;
			{8'd81, 8'd101}: color_data = 12'hf01;
			{8'd81, 8'd102}: color_data = 12'he00;
			{8'd81, 8'd103}: color_data = 12'he00;
			{8'd81, 8'd104}: color_data = 12'he00;
			{8'd81, 8'd105}: color_data = 12'he00;
			{8'd81, 8'd106}: color_data = 12'hc00;
			{8'd81, 8'd117}: color_data = 12'he00;
			{8'd81, 8'd118}: color_data = 12'he00;
			{8'd81, 8'd119}: color_data = 12'he00;
			{8'd81, 8'd120}: color_data = 12'he00;
			{8'd81, 8'd138}: color_data = 12'he00;
			{8'd81, 8'd139}: color_data = 12'he00;
			{8'd81, 8'd140}: color_data = 12'he00;
			{8'd81, 8'd141}: color_data = 12'he00;
			{8'd81, 8'd142}: color_data = 12'he00;
			{8'd81, 8'd143}: color_data = 12'he01;
			{8'd81, 8'd144}: color_data = 12'he00;
			{8'd82, 8'd3}: color_data = 12'h000;
			{8'd82, 8'd4}: color_data = 12'h000;
			{8'd82, 8'd5}: color_data = 12'h100;
			{8'd82, 8'd6}: color_data = 12'hd20;
			{8'd82, 8'd7}: color_data = 12'he21;
			{8'd82, 8'd8}: color_data = 12'he21;
			{8'd82, 8'd9}: color_data = 12'he21;
			{8'd82, 8'd10}: color_data = 12'he21;
			{8'd82, 8'd11}: color_data = 12'he21;
			{8'd82, 8'd12}: color_data = 12'he21;
			{8'd82, 8'd13}: color_data = 12'he21;
			{8'd82, 8'd14}: color_data = 12'he21;
			{8'd82, 8'd15}: color_data = 12'he21;
			{8'd82, 8'd16}: color_data = 12'he21;
			{8'd82, 8'd17}: color_data = 12'he21;
			{8'd82, 8'd18}: color_data = 12'he21;
			{8'd82, 8'd19}: color_data = 12'he21;
			{8'd82, 8'd20}: color_data = 12'he21;
			{8'd82, 8'd21}: color_data = 12'he21;
			{8'd82, 8'd22}: color_data = 12'he21;
			{8'd82, 8'd23}: color_data = 12'he21;
			{8'd82, 8'd24}: color_data = 12'he21;
			{8'd82, 8'd25}: color_data = 12'he21;
			{8'd82, 8'd26}: color_data = 12'he21;
			{8'd82, 8'd27}: color_data = 12'he21;
			{8'd82, 8'd28}: color_data = 12'he21;
			{8'd82, 8'd29}: color_data = 12'hf21;
			{8'd82, 8'd30}: color_data = 12'h810;
			{8'd82, 8'd31}: color_data = 12'h000;
			{8'd82, 8'd32}: color_data = 12'h000;
			{8'd82, 8'd33}: color_data = 12'h000;
			{8'd82, 8'd34}: color_data = 12'h000;
			{8'd82, 8'd35}: color_data = 12'ha80;
			{8'd82, 8'd36}: color_data = 12'hfd0;
			{8'd82, 8'd37}: color_data = 12'hfc0;
			{8'd82, 8'd38}: color_data = 12'hfc0;
			{8'd82, 8'd39}: color_data = 12'hfc0;
			{8'd82, 8'd40}: color_data = 12'hfc0;
			{8'd82, 8'd41}: color_data = 12'hfc0;
			{8'd82, 8'd42}: color_data = 12'hfc0;
			{8'd82, 8'd43}: color_data = 12'hfc0;
			{8'd82, 8'd44}: color_data = 12'hfc0;
			{8'd82, 8'd45}: color_data = 12'hfc0;
			{8'd82, 8'd46}: color_data = 12'hfd0;
			{8'd82, 8'd47}: color_data = 12'hfd0;
			{8'd82, 8'd48}: color_data = 12'hfd0;
			{8'd82, 8'd49}: color_data = 12'hfd0;
			{8'd82, 8'd50}: color_data = 12'hfd0;
			{8'd82, 8'd51}: color_data = 12'hfd0;
			{8'd82, 8'd52}: color_data = 12'hfd0;
			{8'd82, 8'd53}: color_data = 12'hfd0;
			{8'd82, 8'd54}: color_data = 12'hfd0;
			{8'd82, 8'd55}: color_data = 12'hfd0;
			{8'd82, 8'd56}: color_data = 12'hec0;
			{8'd82, 8'd57}: color_data = 12'ha90;
			{8'd82, 8'd58}: color_data = 12'h540;
			{8'd82, 8'd59}: color_data = 12'h110;
			{8'd82, 8'd60}: color_data = 12'h000;
			{8'd82, 8'd61}: color_data = 12'h000;
			{8'd82, 8'd62}: color_data = 12'h000;
			{8'd82, 8'd63}: color_data = 12'h000;
			{8'd82, 8'd64}: color_data = 12'h000;
			{8'd82, 8'd65}: color_data = 12'h120;
			{8'd82, 8'd66}: color_data = 12'h000;
			{8'd82, 8'd67}: color_data = 12'h000;
			{8'd82, 8'd68}: color_data = 12'h000;
			{8'd82, 8'd69}: color_data = 12'h000;
			{8'd82, 8'd70}: color_data = 12'h000;
			{8'd82, 8'd71}: color_data = 12'h000;
			{8'd82, 8'd72}: color_data = 12'h000;
			{8'd82, 8'd73}: color_data = 12'h000;
			{8'd82, 8'd74}: color_data = 12'h000;
			{8'd82, 8'd75}: color_data = 12'h000;
			{8'd82, 8'd100}: color_data = 12'he00;
			{8'd82, 8'd101}: color_data = 12'hf01;
			{8'd82, 8'd102}: color_data = 12'he00;
			{8'd82, 8'd103}: color_data = 12'he00;
			{8'd82, 8'd104}: color_data = 12'he00;
			{8'd82, 8'd105}: color_data = 12'he00;
			{8'd82, 8'd106}: color_data = 12'hc00;
			{8'd82, 8'd117}: color_data = 12'hd01;
			{8'd82, 8'd118}: color_data = 12'he00;
			{8'd82, 8'd138}: color_data = 12'he00;
			{8'd82, 8'd139}: color_data = 12'he00;
			{8'd82, 8'd140}: color_data = 12'he00;
			{8'd82, 8'd141}: color_data = 12'he00;
			{8'd82, 8'd142}: color_data = 12'he00;
			{8'd82, 8'd143}: color_data = 12'he01;
			{8'd82, 8'd144}: color_data = 12'he00;
			{8'd83, 8'd3}: color_data = 12'h000;
			{8'd83, 8'd4}: color_data = 12'h000;
			{8'd83, 8'd5}: color_data = 12'h400;
			{8'd83, 8'd6}: color_data = 12'he21;
			{8'd83, 8'd7}: color_data = 12'he21;
			{8'd83, 8'd8}: color_data = 12'he21;
			{8'd83, 8'd9}: color_data = 12'he21;
			{8'd83, 8'd10}: color_data = 12'he21;
			{8'd83, 8'd11}: color_data = 12'he21;
			{8'd83, 8'd12}: color_data = 12'he21;
			{8'd83, 8'd13}: color_data = 12'he21;
			{8'd83, 8'd14}: color_data = 12'he21;
			{8'd83, 8'd15}: color_data = 12'he21;
			{8'd83, 8'd16}: color_data = 12'he21;
			{8'd83, 8'd17}: color_data = 12'he21;
			{8'd83, 8'd18}: color_data = 12'he21;
			{8'd83, 8'd19}: color_data = 12'he21;
			{8'd83, 8'd20}: color_data = 12'he21;
			{8'd83, 8'd21}: color_data = 12'he21;
			{8'd83, 8'd22}: color_data = 12'he21;
			{8'd83, 8'd23}: color_data = 12'he21;
			{8'd83, 8'd24}: color_data = 12'he21;
			{8'd83, 8'd25}: color_data = 12'he21;
			{8'd83, 8'd26}: color_data = 12'he21;
			{8'd83, 8'd27}: color_data = 12'he21;
			{8'd83, 8'd28}: color_data = 12'he21;
			{8'd83, 8'd29}: color_data = 12'he21;
			{8'd83, 8'd30}: color_data = 12'h710;
			{8'd83, 8'd31}: color_data = 12'h000;
			{8'd83, 8'd32}: color_data = 12'h000;
			{8'd83, 8'd33}: color_data = 12'h000;
			{8'd83, 8'd34}: color_data = 12'h000;
			{8'd83, 8'd35}: color_data = 12'hca0;
			{8'd83, 8'd36}: color_data = 12'hfd0;
			{8'd83, 8'd37}: color_data = 12'hfc0;
			{8'd83, 8'd38}: color_data = 12'hfc0;
			{8'd83, 8'd39}: color_data = 12'hfc0;
			{8'd83, 8'd40}: color_data = 12'hfc0;
			{8'd83, 8'd41}: color_data = 12'hfc0;
			{8'd83, 8'd42}: color_data = 12'hfc0;
			{8'd83, 8'd43}: color_data = 12'hfc0;
			{8'd83, 8'd44}: color_data = 12'hfc0;
			{8'd83, 8'd45}: color_data = 12'hfc0;
			{8'd83, 8'd46}: color_data = 12'hfc0;
			{8'd83, 8'd47}: color_data = 12'hfc0;
			{8'd83, 8'd48}: color_data = 12'hfc0;
			{8'd83, 8'd49}: color_data = 12'hfc0;
			{8'd83, 8'd50}: color_data = 12'hfc0;
			{8'd83, 8'd51}: color_data = 12'hfc0;
			{8'd83, 8'd52}: color_data = 12'hfc0;
			{8'd83, 8'd53}: color_data = 12'hfc0;
			{8'd83, 8'd54}: color_data = 12'hfc0;
			{8'd83, 8'd55}: color_data = 12'hfd0;
			{8'd83, 8'd56}: color_data = 12'hfd0;
			{8'd83, 8'd57}: color_data = 12'hfd0;
			{8'd83, 8'd58}: color_data = 12'hfd0;
			{8'd83, 8'd59}: color_data = 12'heb0;
			{8'd83, 8'd60}: color_data = 12'ha80;
			{8'd83, 8'd61}: color_data = 12'h540;
			{8'd83, 8'd62}: color_data = 12'h100;
			{8'd83, 8'd63}: color_data = 12'h000;
			{8'd83, 8'd64}: color_data = 12'h000;
			{8'd83, 8'd65}: color_data = 12'h000;
			{8'd83, 8'd66}: color_data = 12'h000;
			{8'd83, 8'd67}: color_data = 12'h000;
			{8'd83, 8'd68}: color_data = 12'h000;
			{8'd83, 8'd69}: color_data = 12'h000;
			{8'd83, 8'd70}: color_data = 12'h000;
			{8'd83, 8'd71}: color_data = 12'h000;
			{8'd83, 8'd72}: color_data = 12'h000;
			{8'd83, 8'd73}: color_data = 12'h000;
			{8'd83, 8'd74}: color_data = 12'h000;
			{8'd83, 8'd75}: color_data = 12'h000;
			{8'd83, 8'd100}: color_data = 12'he00;
			{8'd83, 8'd101}: color_data = 12'hf01;
			{8'd83, 8'd102}: color_data = 12'he00;
			{8'd83, 8'd103}: color_data = 12'he00;
			{8'd83, 8'd104}: color_data = 12'he00;
			{8'd83, 8'd105}: color_data = 12'he00;
			{8'd83, 8'd106}: color_data = 12'hc00;
			{8'd83, 8'd121}: color_data = 12'he01;
			{8'd83, 8'd122}: color_data = 12'he00;
			{8'd83, 8'd126}: color_data = 12'hf00;
			{8'd83, 8'd127}: color_data = 12'he00;
			{8'd83, 8'd128}: color_data = 12'he00;
			{8'd83, 8'd129}: color_data = 12'he00;
			{8'd83, 8'd130}: color_data = 12'he00;
			{8'd83, 8'd131}: color_data = 12'he00;
			{8'd83, 8'd138}: color_data = 12'he00;
			{8'd83, 8'd139}: color_data = 12'he00;
			{8'd83, 8'd140}: color_data = 12'he00;
			{8'd83, 8'd141}: color_data = 12'he00;
			{8'd83, 8'd142}: color_data = 12'he00;
			{8'd83, 8'd143}: color_data = 12'he01;
			{8'd83, 8'd144}: color_data = 12'he00;
			{8'd84, 8'd3}: color_data = 12'h000;
			{8'd84, 8'd4}: color_data = 12'h000;
			{8'd84, 8'd5}: color_data = 12'h610;
			{8'd84, 8'd6}: color_data = 12'he21;
			{8'd84, 8'd7}: color_data = 12'he21;
			{8'd84, 8'd8}: color_data = 12'he21;
			{8'd84, 8'd9}: color_data = 12'he21;
			{8'd84, 8'd10}: color_data = 12'he21;
			{8'd84, 8'd11}: color_data = 12'he21;
			{8'd84, 8'd12}: color_data = 12'he21;
			{8'd84, 8'd13}: color_data = 12'he21;
			{8'd84, 8'd14}: color_data = 12'he21;
			{8'd84, 8'd15}: color_data = 12'he21;
			{8'd84, 8'd16}: color_data = 12'he21;
			{8'd84, 8'd17}: color_data = 12'he21;
			{8'd84, 8'd18}: color_data = 12'he21;
			{8'd84, 8'd19}: color_data = 12'he21;
			{8'd84, 8'd20}: color_data = 12'he21;
			{8'd84, 8'd21}: color_data = 12'he21;
			{8'd84, 8'd22}: color_data = 12'he21;
			{8'd84, 8'd23}: color_data = 12'he21;
			{8'd84, 8'd24}: color_data = 12'he21;
			{8'd84, 8'd25}: color_data = 12'he21;
			{8'd84, 8'd26}: color_data = 12'he21;
			{8'd84, 8'd27}: color_data = 12'he21;
			{8'd84, 8'd28}: color_data = 12'he21;
			{8'd84, 8'd29}: color_data = 12'he21;
			{8'd84, 8'd30}: color_data = 12'h500;
			{8'd84, 8'd31}: color_data = 12'h000;
			{8'd84, 8'd32}: color_data = 12'h000;
			{8'd84, 8'd33}: color_data = 12'h000;
			{8'd84, 8'd34}: color_data = 12'h110;
			{8'd84, 8'd35}: color_data = 12'heb0;
			{8'd84, 8'd36}: color_data = 12'hfd0;
			{8'd84, 8'd37}: color_data = 12'hfc0;
			{8'd84, 8'd38}: color_data = 12'hfc0;
			{8'd84, 8'd39}: color_data = 12'hfc0;
			{8'd84, 8'd40}: color_data = 12'hfc0;
			{8'd84, 8'd41}: color_data = 12'hfc0;
			{8'd84, 8'd42}: color_data = 12'hfc0;
			{8'd84, 8'd43}: color_data = 12'hfc0;
			{8'd84, 8'd44}: color_data = 12'hfc0;
			{8'd84, 8'd45}: color_data = 12'hfc0;
			{8'd84, 8'd46}: color_data = 12'hfc0;
			{8'd84, 8'd47}: color_data = 12'hfc0;
			{8'd84, 8'd48}: color_data = 12'hfc0;
			{8'd84, 8'd49}: color_data = 12'hfc0;
			{8'd84, 8'd50}: color_data = 12'hfc0;
			{8'd84, 8'd51}: color_data = 12'hfc0;
			{8'd84, 8'd52}: color_data = 12'hfc0;
			{8'd84, 8'd53}: color_data = 12'hfc0;
			{8'd84, 8'd54}: color_data = 12'hfc0;
			{8'd84, 8'd55}: color_data = 12'hfc0;
			{8'd84, 8'd56}: color_data = 12'hfc0;
			{8'd84, 8'd57}: color_data = 12'hfc0;
			{8'd84, 8'd58}: color_data = 12'hfc0;
			{8'd84, 8'd59}: color_data = 12'hfd0;
			{8'd84, 8'd60}: color_data = 12'hfd0;
			{8'd84, 8'd61}: color_data = 12'hfd0;
			{8'd84, 8'd62}: color_data = 12'heb0;
			{8'd84, 8'd63}: color_data = 12'h970;
			{8'd84, 8'd64}: color_data = 12'h430;
			{8'd84, 8'd65}: color_data = 12'h000;
			{8'd84, 8'd66}: color_data = 12'h000;
			{8'd84, 8'd67}: color_data = 12'h000;
			{8'd84, 8'd68}: color_data = 12'h000;
			{8'd84, 8'd69}: color_data = 12'h000;
			{8'd84, 8'd70}: color_data = 12'h000;
			{8'd84, 8'd71}: color_data = 12'h000;
			{8'd84, 8'd72}: color_data = 12'h000;
			{8'd84, 8'd73}: color_data = 12'h000;
			{8'd84, 8'd74}: color_data = 12'h000;
			{8'd84, 8'd75}: color_data = 12'h000;
			{8'd84, 8'd100}: color_data = 12'he00;
			{8'd84, 8'd101}: color_data = 12'hf01;
			{8'd84, 8'd102}: color_data = 12'he00;
			{8'd84, 8'd103}: color_data = 12'he00;
			{8'd84, 8'd104}: color_data = 12'he00;
			{8'd84, 8'd105}: color_data = 12'he00;
			{8'd84, 8'd106}: color_data = 12'hc00;
			{8'd84, 8'd119}: color_data = 12'he00;
			{8'd84, 8'd120}: color_data = 12'he00;
			{8'd84, 8'd121}: color_data = 12'he00;
			{8'd84, 8'd122}: color_data = 12'he00;
			{8'd84, 8'd125}: color_data = 12'hc00;
			{8'd84, 8'd126}: color_data = 12'he00;
			{8'd84, 8'd127}: color_data = 12'he01;
			{8'd84, 8'd128}: color_data = 12'he01;
			{8'd84, 8'd129}: color_data = 12'he01;
			{8'd84, 8'd130}: color_data = 12'hf01;
			{8'd84, 8'd131}: color_data = 12'he00;
			{8'd84, 8'd132}: color_data = 12'he00;
			{8'd84, 8'd138}: color_data = 12'he00;
			{8'd84, 8'd139}: color_data = 12'he00;
			{8'd84, 8'd140}: color_data = 12'he00;
			{8'd84, 8'd141}: color_data = 12'he00;
			{8'd84, 8'd142}: color_data = 12'he00;
			{8'd84, 8'd143}: color_data = 12'he01;
			{8'd84, 8'd144}: color_data = 12'he00;
			{8'd85, 8'd2}: color_data = 12'h000;
			{8'd85, 8'd3}: color_data = 12'h000;
			{8'd85, 8'd4}: color_data = 12'h000;
			{8'd85, 8'd5}: color_data = 12'h910;
			{8'd85, 8'd6}: color_data = 12'he21;
			{8'd85, 8'd7}: color_data = 12'he21;
			{8'd85, 8'd8}: color_data = 12'he21;
			{8'd85, 8'd9}: color_data = 12'he21;
			{8'd85, 8'd10}: color_data = 12'he21;
			{8'd85, 8'd11}: color_data = 12'he21;
			{8'd85, 8'd12}: color_data = 12'he21;
			{8'd85, 8'd13}: color_data = 12'he21;
			{8'd85, 8'd14}: color_data = 12'he21;
			{8'd85, 8'd15}: color_data = 12'he21;
			{8'd85, 8'd16}: color_data = 12'he21;
			{8'd85, 8'd17}: color_data = 12'he21;
			{8'd85, 8'd18}: color_data = 12'he21;
			{8'd85, 8'd19}: color_data = 12'he21;
			{8'd85, 8'd20}: color_data = 12'he21;
			{8'd85, 8'd21}: color_data = 12'he21;
			{8'd85, 8'd22}: color_data = 12'he21;
			{8'd85, 8'd23}: color_data = 12'he21;
			{8'd85, 8'd24}: color_data = 12'he21;
			{8'd85, 8'd25}: color_data = 12'he21;
			{8'd85, 8'd26}: color_data = 12'he21;
			{8'd85, 8'd27}: color_data = 12'he21;
			{8'd85, 8'd28}: color_data = 12'he21;
			{8'd85, 8'd29}: color_data = 12'he21;
			{8'd85, 8'd30}: color_data = 12'h400;
			{8'd85, 8'd31}: color_data = 12'h000;
			{8'd85, 8'd32}: color_data = 12'h000;
			{8'd85, 8'd33}: color_data = 12'h000;
			{8'd85, 8'd34}: color_data = 12'h220;
			{8'd85, 8'd35}: color_data = 12'hfc0;
			{8'd85, 8'd36}: color_data = 12'hfd0;
			{8'd85, 8'd37}: color_data = 12'hfc0;
			{8'd85, 8'd38}: color_data = 12'hfc0;
			{8'd85, 8'd39}: color_data = 12'hfc0;
			{8'd85, 8'd40}: color_data = 12'hfc0;
			{8'd85, 8'd41}: color_data = 12'hfc0;
			{8'd85, 8'd42}: color_data = 12'hfc0;
			{8'd85, 8'd43}: color_data = 12'hfc0;
			{8'd85, 8'd44}: color_data = 12'hfc0;
			{8'd85, 8'd45}: color_data = 12'hfc0;
			{8'd85, 8'd46}: color_data = 12'hfc0;
			{8'd85, 8'd47}: color_data = 12'hfc0;
			{8'd85, 8'd48}: color_data = 12'hfc0;
			{8'd85, 8'd49}: color_data = 12'hfc0;
			{8'd85, 8'd50}: color_data = 12'hfc0;
			{8'd85, 8'd51}: color_data = 12'hfc0;
			{8'd85, 8'd52}: color_data = 12'hfc0;
			{8'd85, 8'd53}: color_data = 12'hfc0;
			{8'd85, 8'd54}: color_data = 12'hfc0;
			{8'd85, 8'd55}: color_data = 12'hfc0;
			{8'd85, 8'd56}: color_data = 12'hfc0;
			{8'd85, 8'd57}: color_data = 12'hfc0;
			{8'd85, 8'd58}: color_data = 12'hfc0;
			{8'd85, 8'd59}: color_data = 12'hfc0;
			{8'd85, 8'd60}: color_data = 12'hfc0;
			{8'd85, 8'd61}: color_data = 12'hfc0;
			{8'd85, 8'd62}: color_data = 12'hfd0;
			{8'd85, 8'd63}: color_data = 12'hfd0;
			{8'd85, 8'd64}: color_data = 12'hfd0;
			{8'd85, 8'd65}: color_data = 12'hdb0;
			{8'd85, 8'd66}: color_data = 12'h870;
			{8'd85, 8'd67}: color_data = 12'h320;
			{8'd85, 8'd68}: color_data = 12'h000;
			{8'd85, 8'd69}: color_data = 12'h000;
			{8'd85, 8'd70}: color_data = 12'h000;
			{8'd85, 8'd71}: color_data = 12'h000;
			{8'd85, 8'd72}: color_data = 12'h000;
			{8'd85, 8'd73}: color_data = 12'h000;
			{8'd85, 8'd74}: color_data = 12'h000;
			{8'd85, 8'd100}: color_data = 12'he00;
			{8'd85, 8'd101}: color_data = 12'hf01;
			{8'd85, 8'd102}: color_data = 12'he00;
			{8'd85, 8'd103}: color_data = 12'he00;
			{8'd85, 8'd104}: color_data = 12'he00;
			{8'd85, 8'd105}: color_data = 12'he00;
			{8'd85, 8'd106}: color_data = 12'hc00;
			{8'd85, 8'd118}: color_data = 12'hd00;
			{8'd85, 8'd119}: color_data = 12'he00;
			{8'd85, 8'd120}: color_data = 12'hf01;
			{8'd85, 8'd121}: color_data = 12'hf01;
			{8'd85, 8'd122}: color_data = 12'he00;
			{8'd85, 8'd125}: color_data = 12'he00;
			{8'd85, 8'd126}: color_data = 12'hf01;
			{8'd85, 8'd127}: color_data = 12'he00;
			{8'd85, 8'd128}: color_data = 12'he00;
			{8'd85, 8'd129}: color_data = 12'he00;
			{8'd85, 8'd130}: color_data = 12'he00;
			{8'd85, 8'd131}: color_data = 12'he00;
			{8'd85, 8'd132}: color_data = 12'he00;
			{8'd85, 8'd133}: color_data = 12'hd00;
			{8'd85, 8'd138}: color_data = 12'he00;
			{8'd85, 8'd139}: color_data = 12'he00;
			{8'd85, 8'd140}: color_data = 12'he00;
			{8'd85, 8'd141}: color_data = 12'he00;
			{8'd85, 8'd142}: color_data = 12'he00;
			{8'd85, 8'd143}: color_data = 12'he01;
			{8'd85, 8'd144}: color_data = 12'he00;
			{8'd86, 8'd2}: color_data = 12'h000;
			{8'd86, 8'd3}: color_data = 12'h000;
			{8'd86, 8'd4}: color_data = 12'h000;
			{8'd86, 8'd5}: color_data = 12'hb10;
			{8'd86, 8'd6}: color_data = 12'he21;
			{8'd86, 8'd7}: color_data = 12'he21;
			{8'd86, 8'd8}: color_data = 12'he21;
			{8'd86, 8'd9}: color_data = 12'he21;
			{8'd86, 8'd10}: color_data = 12'he21;
			{8'd86, 8'd11}: color_data = 12'he21;
			{8'd86, 8'd12}: color_data = 12'he21;
			{8'd86, 8'd13}: color_data = 12'he21;
			{8'd86, 8'd14}: color_data = 12'he21;
			{8'd86, 8'd15}: color_data = 12'he21;
			{8'd86, 8'd16}: color_data = 12'he21;
			{8'd86, 8'd17}: color_data = 12'he21;
			{8'd86, 8'd18}: color_data = 12'he21;
			{8'd86, 8'd19}: color_data = 12'he21;
			{8'd86, 8'd20}: color_data = 12'he21;
			{8'd86, 8'd21}: color_data = 12'he21;
			{8'd86, 8'd22}: color_data = 12'he21;
			{8'd86, 8'd23}: color_data = 12'he21;
			{8'd86, 8'd24}: color_data = 12'he21;
			{8'd86, 8'd25}: color_data = 12'he21;
			{8'd86, 8'd26}: color_data = 12'he21;
			{8'd86, 8'd27}: color_data = 12'he21;
			{8'd86, 8'd28}: color_data = 12'he21;
			{8'd86, 8'd29}: color_data = 12'he21;
			{8'd86, 8'd30}: color_data = 12'h300;
			{8'd86, 8'd31}: color_data = 12'h000;
			{8'd86, 8'd32}: color_data = 12'h000;
			{8'd86, 8'd33}: color_data = 12'h000;
			{8'd86, 8'd34}: color_data = 12'h540;
			{8'd86, 8'd35}: color_data = 12'hfd0;
			{8'd86, 8'd36}: color_data = 12'hfc0;
			{8'd86, 8'd37}: color_data = 12'hfc0;
			{8'd86, 8'd38}: color_data = 12'hfc0;
			{8'd86, 8'd39}: color_data = 12'hfc0;
			{8'd86, 8'd40}: color_data = 12'hfc0;
			{8'd86, 8'd41}: color_data = 12'hfc0;
			{8'd86, 8'd42}: color_data = 12'hfc0;
			{8'd86, 8'd43}: color_data = 12'hfc0;
			{8'd86, 8'd44}: color_data = 12'hfc0;
			{8'd86, 8'd45}: color_data = 12'hfc0;
			{8'd86, 8'd46}: color_data = 12'hfc0;
			{8'd86, 8'd47}: color_data = 12'hfc0;
			{8'd86, 8'd48}: color_data = 12'hfc0;
			{8'd86, 8'd49}: color_data = 12'hfc0;
			{8'd86, 8'd50}: color_data = 12'hfc0;
			{8'd86, 8'd51}: color_data = 12'hfc0;
			{8'd86, 8'd52}: color_data = 12'hfc0;
			{8'd86, 8'd53}: color_data = 12'hfc0;
			{8'd86, 8'd54}: color_data = 12'hfc0;
			{8'd86, 8'd55}: color_data = 12'hfc0;
			{8'd86, 8'd56}: color_data = 12'hfc0;
			{8'd86, 8'd57}: color_data = 12'hfc0;
			{8'd86, 8'd58}: color_data = 12'hfc0;
			{8'd86, 8'd59}: color_data = 12'hfc0;
			{8'd86, 8'd60}: color_data = 12'hfc0;
			{8'd86, 8'd61}: color_data = 12'hfc0;
			{8'd86, 8'd62}: color_data = 12'hfc0;
			{8'd86, 8'd63}: color_data = 12'hfc0;
			{8'd86, 8'd64}: color_data = 12'hfc0;
			{8'd86, 8'd65}: color_data = 12'hfd0;
			{8'd86, 8'd66}: color_data = 12'hfd0;
			{8'd86, 8'd67}: color_data = 12'hdb0;
			{8'd86, 8'd68}: color_data = 12'h000;
			{8'd86, 8'd69}: color_data = 12'h000;
			{8'd86, 8'd70}: color_data = 12'h000;
			{8'd86, 8'd71}: color_data = 12'h000;
			{8'd86, 8'd72}: color_data = 12'h000;
			{8'd86, 8'd73}: color_data = 12'h000;
			{8'd86, 8'd74}: color_data = 12'h000;
			{8'd86, 8'd100}: color_data = 12'he00;
			{8'd86, 8'd101}: color_data = 12'hf01;
			{8'd86, 8'd102}: color_data = 12'he00;
			{8'd86, 8'd103}: color_data = 12'he00;
			{8'd86, 8'd104}: color_data = 12'he00;
			{8'd86, 8'd105}: color_data = 12'he00;
			{8'd86, 8'd106}: color_data = 12'hc00;
			{8'd86, 8'd118}: color_data = 12'he00;
			{8'd86, 8'd119}: color_data = 12'hf01;
			{8'd86, 8'd120}: color_data = 12'he00;
			{8'd86, 8'd121}: color_data = 12'he01;
			{8'd86, 8'd122}: color_data = 12'he00;
			{8'd86, 8'd124}: color_data = 12'hf00;
			{8'd86, 8'd125}: color_data = 12'he00;
			{8'd86, 8'd126}: color_data = 12'he00;
			{8'd86, 8'd127}: color_data = 12'he00;
			{8'd86, 8'd128}: color_data = 12'he00;
			{8'd86, 8'd129}: color_data = 12'he00;
			{8'd86, 8'd130}: color_data = 12'he00;
			{8'd86, 8'd131}: color_data = 12'he00;
			{8'd86, 8'd132}: color_data = 12'hf01;
			{8'd86, 8'd133}: color_data = 12'he00;
			{8'd86, 8'd138}: color_data = 12'he00;
			{8'd86, 8'd139}: color_data = 12'he00;
			{8'd86, 8'd140}: color_data = 12'he00;
			{8'd86, 8'd141}: color_data = 12'he00;
			{8'd86, 8'd142}: color_data = 12'he00;
			{8'd86, 8'd143}: color_data = 12'he01;
			{8'd86, 8'd144}: color_data = 12'he00;
			{8'd87, 8'd2}: color_data = 12'h000;
			{8'd87, 8'd3}: color_data = 12'h000;
			{8'd87, 8'd4}: color_data = 12'h100;
			{8'd87, 8'd5}: color_data = 12'hd20;
			{8'd87, 8'd6}: color_data = 12'he21;
			{8'd87, 8'd7}: color_data = 12'he21;
			{8'd87, 8'd8}: color_data = 12'he21;
			{8'd87, 8'd9}: color_data = 12'he21;
			{8'd87, 8'd10}: color_data = 12'h810;
			{8'd87, 8'd11}: color_data = 12'h200;
			{8'd87, 8'd12}: color_data = 12'h300;
			{8'd87, 8'd13}: color_data = 12'h400;
			{8'd87, 8'd14}: color_data = 12'h500;
			{8'd87, 8'd15}: color_data = 12'h600;
			{8'd87, 8'd16}: color_data = 12'h710;
			{8'd87, 8'd17}: color_data = 12'h710;
			{8'd87, 8'd18}: color_data = 12'hc10;
			{8'd87, 8'd19}: color_data = 12'he21;
			{8'd87, 8'd20}: color_data = 12'he21;
			{8'd87, 8'd21}: color_data = 12'he21;
			{8'd87, 8'd22}: color_data = 12'he21;
			{8'd87, 8'd23}: color_data = 12'hd20;
			{8'd87, 8'd24}: color_data = 12'hc20;
			{8'd87, 8'd25}: color_data = 12'hd20;
			{8'd87, 8'd26}: color_data = 12'hd20;
			{8'd87, 8'd27}: color_data = 12'he21;
			{8'd87, 8'd28}: color_data = 12'he21;
			{8'd87, 8'd29}: color_data = 12'he20;
			{8'd87, 8'd30}: color_data = 12'h200;
			{8'd87, 8'd31}: color_data = 12'h000;
			{8'd87, 8'd32}: color_data = 12'h000;
			{8'd87, 8'd33}: color_data = 12'h000;
			{8'd87, 8'd34}: color_data = 12'h760;
			{8'd87, 8'd35}: color_data = 12'hfd0;
			{8'd87, 8'd36}: color_data = 12'hfc0;
			{8'd87, 8'd37}: color_data = 12'hfc0;
			{8'd87, 8'd38}: color_data = 12'hfc0;
			{8'd87, 8'd39}: color_data = 12'hfc0;
			{8'd87, 8'd40}: color_data = 12'hfc0;
			{8'd87, 8'd41}: color_data = 12'hfc0;
			{8'd87, 8'd42}: color_data = 12'hfc0;
			{8'd87, 8'd43}: color_data = 12'hfc0;
			{8'd87, 8'd44}: color_data = 12'hfc0;
			{8'd87, 8'd45}: color_data = 12'hfc0;
			{8'd87, 8'd46}: color_data = 12'hfc0;
			{8'd87, 8'd47}: color_data = 12'hfc0;
			{8'd87, 8'd48}: color_data = 12'hfc0;
			{8'd87, 8'd49}: color_data = 12'hfc0;
			{8'd87, 8'd50}: color_data = 12'hfc0;
			{8'd87, 8'd51}: color_data = 12'hfc0;
			{8'd87, 8'd52}: color_data = 12'hfc0;
			{8'd87, 8'd53}: color_data = 12'hfc0;
			{8'd87, 8'd54}: color_data = 12'hfc0;
			{8'd87, 8'd55}: color_data = 12'hfc0;
			{8'd87, 8'd56}: color_data = 12'hfc0;
			{8'd87, 8'd57}: color_data = 12'hfc0;
			{8'd87, 8'd58}: color_data = 12'hfc0;
			{8'd87, 8'd59}: color_data = 12'hfc0;
			{8'd87, 8'd60}: color_data = 12'hfc0;
			{8'd87, 8'd61}: color_data = 12'hfc0;
			{8'd87, 8'd62}: color_data = 12'hfc0;
			{8'd87, 8'd63}: color_data = 12'hfc0;
			{8'd87, 8'd64}: color_data = 12'hfc0;
			{8'd87, 8'd65}: color_data = 12'hfc0;
			{8'd87, 8'd66}: color_data = 12'hfd0;
			{8'd87, 8'd67}: color_data = 12'hca0;
			{8'd87, 8'd68}: color_data = 12'h000;
			{8'd87, 8'd69}: color_data = 12'h000;
			{8'd87, 8'd70}: color_data = 12'h000;
			{8'd87, 8'd71}: color_data = 12'h000;
			{8'd87, 8'd72}: color_data = 12'h000;
			{8'd87, 8'd73}: color_data = 12'h000;
			{8'd87, 8'd74}: color_data = 12'h000;
			{8'd87, 8'd100}: color_data = 12'he00;
			{8'd87, 8'd101}: color_data = 12'hf01;
			{8'd87, 8'd102}: color_data = 12'he00;
			{8'd87, 8'd103}: color_data = 12'he00;
			{8'd87, 8'd104}: color_data = 12'he00;
			{8'd87, 8'd105}: color_data = 12'he00;
			{8'd87, 8'd106}: color_data = 12'hc00;
			{8'd87, 8'd117}: color_data = 12'he00;
			{8'd87, 8'd118}: color_data = 12'he00;
			{8'd87, 8'd119}: color_data = 12'he00;
			{8'd87, 8'd120}: color_data = 12'he00;
			{8'd87, 8'd121}: color_data = 12'he00;
			{8'd87, 8'd122}: color_data = 12'he00;
			{8'd87, 8'd124}: color_data = 12'he00;
			{8'd87, 8'd125}: color_data = 12'he00;
			{8'd87, 8'd126}: color_data = 12'he00;
			{8'd87, 8'd127}: color_data = 12'he00;
			{8'd87, 8'd128}: color_data = 12'he00;
			{8'd87, 8'd129}: color_data = 12'he00;
			{8'd87, 8'd130}: color_data = 12'he00;
			{8'd87, 8'd131}: color_data = 12'he00;
			{8'd87, 8'd132}: color_data = 12'he00;
			{8'd87, 8'd133}: color_data = 12'he00;
			{8'd87, 8'd138}: color_data = 12'he00;
			{8'd87, 8'd139}: color_data = 12'he00;
			{8'd87, 8'd140}: color_data = 12'he00;
			{8'd87, 8'd141}: color_data = 12'he00;
			{8'd87, 8'd142}: color_data = 12'he00;
			{8'd87, 8'd143}: color_data = 12'he01;
			{8'd87, 8'd144}: color_data = 12'he00;
			{8'd88, 8'd2}: color_data = 12'h000;
			{8'd88, 8'd3}: color_data = 12'h000;
			{8'd88, 8'd4}: color_data = 12'h300;
			{8'd88, 8'd5}: color_data = 12'he21;
			{8'd88, 8'd6}: color_data = 12'he21;
			{8'd88, 8'd7}: color_data = 12'he21;
			{8'd88, 8'd8}: color_data = 12'he21;
			{8'd88, 8'd9}: color_data = 12'he21;
			{8'd88, 8'd10}: color_data = 12'hb10;
			{8'd88, 8'd11}: color_data = 12'h000;
			{8'd88, 8'd12}: color_data = 12'h000;
			{8'd88, 8'd13}: color_data = 12'h000;
			{8'd88, 8'd14}: color_data = 12'h000;
			{8'd88, 8'd15}: color_data = 12'h000;
			{8'd88, 8'd16}: color_data = 12'h000;
			{8'd88, 8'd17}: color_data = 12'h000;
			{8'd88, 8'd18}: color_data = 12'hb10;
			{8'd88, 8'd19}: color_data = 12'he21;
			{8'd88, 8'd20}: color_data = 12'he21;
			{8'd88, 8'd21}: color_data = 12'he21;
			{8'd88, 8'd22}: color_data = 12'he21;
			{8'd88, 8'd23}: color_data = 12'ha10;
			{8'd88, 8'd24}: color_data = 12'h000;
			{8'd88, 8'd25}: color_data = 12'h100;
			{8'd88, 8'd26}: color_data = 12'h200;
			{8'd88, 8'd27}: color_data = 12'h200;
			{8'd88, 8'd28}: color_data = 12'h300;
			{8'd88, 8'd29}: color_data = 12'h300;
			{8'd88, 8'd30}: color_data = 12'h000;
			{8'd88, 8'd31}: color_data = 12'h000;
			{8'd88, 8'd32}: color_data = 12'h000;
			{8'd88, 8'd33}: color_data = 12'h000;
			{8'd88, 8'd34}: color_data = 12'h980;
			{8'd88, 8'd35}: color_data = 12'hfd0;
			{8'd88, 8'd36}: color_data = 12'hfc0;
			{8'd88, 8'd37}: color_data = 12'hfc0;
			{8'd88, 8'd38}: color_data = 12'hfc0;
			{8'd88, 8'd39}: color_data = 12'hfc0;
			{8'd88, 8'd40}: color_data = 12'hfc0;
			{8'd88, 8'd41}: color_data = 12'hfc0;
			{8'd88, 8'd42}: color_data = 12'hfc0;
			{8'd88, 8'd43}: color_data = 12'hfc0;
			{8'd88, 8'd44}: color_data = 12'hfc0;
			{8'd88, 8'd45}: color_data = 12'hfc0;
			{8'd88, 8'd46}: color_data = 12'hfc0;
			{8'd88, 8'd47}: color_data = 12'hfc0;
			{8'd88, 8'd48}: color_data = 12'hfc0;
			{8'd88, 8'd49}: color_data = 12'hfc0;
			{8'd88, 8'd50}: color_data = 12'hfc0;
			{8'd88, 8'd51}: color_data = 12'hfc0;
			{8'd88, 8'd52}: color_data = 12'hfc0;
			{8'd88, 8'd53}: color_data = 12'hfc0;
			{8'd88, 8'd54}: color_data = 12'hfc0;
			{8'd88, 8'd55}: color_data = 12'hfc0;
			{8'd88, 8'd56}: color_data = 12'hfc0;
			{8'd88, 8'd57}: color_data = 12'hfc0;
			{8'd88, 8'd58}: color_data = 12'hfc0;
			{8'd88, 8'd59}: color_data = 12'hfc0;
			{8'd88, 8'd60}: color_data = 12'hfc0;
			{8'd88, 8'd61}: color_data = 12'hfc0;
			{8'd88, 8'd62}: color_data = 12'hfc0;
			{8'd88, 8'd63}: color_data = 12'hfc0;
			{8'd88, 8'd64}: color_data = 12'hfc0;
			{8'd88, 8'd65}: color_data = 12'hfc0;
			{8'd88, 8'd66}: color_data = 12'hfd0;
			{8'd88, 8'd67}: color_data = 12'hb90;
			{8'd88, 8'd68}: color_data = 12'h000;
			{8'd88, 8'd69}: color_data = 12'h000;
			{8'd88, 8'd70}: color_data = 12'h000;
			{8'd88, 8'd71}: color_data = 12'h000;
			{8'd88, 8'd72}: color_data = 12'h000;
			{8'd88, 8'd73}: color_data = 12'h000;
			{8'd88, 8'd74}: color_data = 12'h000;
			{8'd88, 8'd100}: color_data = 12'he00;
			{8'd88, 8'd101}: color_data = 12'hf01;
			{8'd88, 8'd102}: color_data = 12'he00;
			{8'd88, 8'd103}: color_data = 12'he00;
			{8'd88, 8'd104}: color_data = 12'he00;
			{8'd88, 8'd105}: color_data = 12'he00;
			{8'd88, 8'd106}: color_data = 12'hc00;
			{8'd88, 8'd117}: color_data = 12'he00;
			{8'd88, 8'd118}: color_data = 12'he00;
			{8'd88, 8'd119}: color_data = 12'he00;
			{8'd88, 8'd120}: color_data = 12'he00;
			{8'd88, 8'd121}: color_data = 12'he00;
			{8'd88, 8'd122}: color_data = 12'he00;
			{8'd88, 8'd124}: color_data = 12'he00;
			{8'd88, 8'd125}: color_data = 12'he00;
			{8'd88, 8'd126}: color_data = 12'he00;
			{8'd88, 8'd127}: color_data = 12'he00;
			{8'd88, 8'd128}: color_data = 12'he00;
			{8'd88, 8'd129}: color_data = 12'he01;
			{8'd88, 8'd130}: color_data = 12'he00;
			{8'd88, 8'd131}: color_data = 12'he00;
			{8'd88, 8'd132}: color_data = 12'he00;
			{8'd88, 8'd133}: color_data = 12'he00;
			{8'd88, 8'd134}: color_data = 12'hf00;
			{8'd88, 8'd138}: color_data = 12'he00;
			{8'd88, 8'd139}: color_data = 12'he00;
			{8'd88, 8'd140}: color_data = 12'he00;
			{8'd88, 8'd141}: color_data = 12'he00;
			{8'd88, 8'd142}: color_data = 12'he00;
			{8'd88, 8'd143}: color_data = 12'he01;
			{8'd88, 8'd144}: color_data = 12'he00;
			{8'd89, 8'd2}: color_data = 12'h000;
			{8'd89, 8'd3}: color_data = 12'h000;
			{8'd89, 8'd4}: color_data = 12'h500;
			{8'd89, 8'd5}: color_data = 12'he21;
			{8'd89, 8'd6}: color_data = 12'he21;
			{8'd89, 8'd7}: color_data = 12'he21;
			{8'd89, 8'd8}: color_data = 12'he21;
			{8'd89, 8'd9}: color_data = 12'he21;
			{8'd89, 8'd10}: color_data = 12'he21;
			{8'd89, 8'd11}: color_data = 12'h300;
			{8'd89, 8'd12}: color_data = 12'h000;
			{8'd89, 8'd13}: color_data = 12'h000;
			{8'd89, 8'd14}: color_data = 12'h000;
			{8'd89, 8'd15}: color_data = 12'h000;
			{8'd89, 8'd16}: color_data = 12'h000;
			{8'd89, 8'd17}: color_data = 12'h100;
			{8'd89, 8'd18}: color_data = 12'hd20;
			{8'd89, 8'd19}: color_data = 12'he21;
			{8'd89, 8'd20}: color_data = 12'he21;
			{8'd89, 8'd21}: color_data = 12'he21;
			{8'd89, 8'd22}: color_data = 12'he21;
			{8'd89, 8'd23}: color_data = 12'h910;
			{8'd89, 8'd24}: color_data = 12'h000;
			{8'd89, 8'd25}: color_data = 12'h000;
			{8'd89, 8'd26}: color_data = 12'h000;
			{8'd89, 8'd27}: color_data = 12'h000;
			{8'd89, 8'd28}: color_data = 12'h000;
			{8'd89, 8'd29}: color_data = 12'h000;
			{8'd89, 8'd30}: color_data = 12'h000;
			{8'd89, 8'd31}: color_data = 12'h000;
			{8'd89, 8'd32}: color_data = 12'h000;
			{8'd89, 8'd33}: color_data = 12'h000;
			{8'd89, 8'd34}: color_data = 12'hca0;
			{8'd89, 8'd35}: color_data = 12'hfd0;
			{8'd89, 8'd36}: color_data = 12'hfc0;
			{8'd89, 8'd37}: color_data = 12'hfc0;
			{8'd89, 8'd38}: color_data = 12'hfc0;
			{8'd89, 8'd39}: color_data = 12'hfc0;
			{8'd89, 8'd40}: color_data = 12'hfc0;
			{8'd89, 8'd41}: color_data = 12'hfc0;
			{8'd89, 8'd42}: color_data = 12'hfc0;
			{8'd89, 8'd43}: color_data = 12'hfc0;
			{8'd89, 8'd44}: color_data = 12'hfc0;
			{8'd89, 8'd45}: color_data = 12'hfc0;
			{8'd89, 8'd46}: color_data = 12'hfc0;
			{8'd89, 8'd47}: color_data = 12'hfc0;
			{8'd89, 8'd48}: color_data = 12'hfc0;
			{8'd89, 8'd49}: color_data = 12'hfc0;
			{8'd89, 8'd50}: color_data = 12'hfc0;
			{8'd89, 8'd51}: color_data = 12'hfc0;
			{8'd89, 8'd52}: color_data = 12'hfc0;
			{8'd89, 8'd53}: color_data = 12'hfc0;
			{8'd89, 8'd54}: color_data = 12'hfc0;
			{8'd89, 8'd55}: color_data = 12'hfc0;
			{8'd89, 8'd56}: color_data = 12'hfc0;
			{8'd89, 8'd57}: color_data = 12'hfc0;
			{8'd89, 8'd58}: color_data = 12'hfc0;
			{8'd89, 8'd59}: color_data = 12'hfc0;
			{8'd89, 8'd60}: color_data = 12'hfc0;
			{8'd89, 8'd61}: color_data = 12'hfc0;
			{8'd89, 8'd62}: color_data = 12'hfc0;
			{8'd89, 8'd63}: color_data = 12'hfc0;
			{8'd89, 8'd64}: color_data = 12'hfc0;
			{8'd89, 8'd65}: color_data = 12'hfc0;
			{8'd89, 8'd66}: color_data = 12'hfd0;
			{8'd89, 8'd67}: color_data = 12'ha80;
			{8'd89, 8'd68}: color_data = 12'h000;
			{8'd89, 8'd69}: color_data = 12'h000;
			{8'd89, 8'd70}: color_data = 12'h000;
			{8'd89, 8'd71}: color_data = 12'h000;
			{8'd89, 8'd72}: color_data = 12'h000;
			{8'd89, 8'd73}: color_data = 12'h000;
			{8'd89, 8'd74}: color_data = 12'h000;
			{8'd89, 8'd100}: color_data = 12'he00;
			{8'd89, 8'd101}: color_data = 12'hf01;
			{8'd89, 8'd102}: color_data = 12'he00;
			{8'd89, 8'd103}: color_data = 12'he00;
			{8'd89, 8'd104}: color_data = 12'he00;
			{8'd89, 8'd105}: color_data = 12'he00;
			{8'd89, 8'd106}: color_data = 12'hc00;
			{8'd89, 8'd117}: color_data = 12'he01;
			{8'd89, 8'd118}: color_data = 12'he01;
			{8'd89, 8'd119}: color_data = 12'he00;
			{8'd89, 8'd120}: color_data = 12'he00;
			{8'd89, 8'd121}: color_data = 12'he00;
			{8'd89, 8'd122}: color_data = 12'he00;
			{8'd89, 8'd124}: color_data = 12'he00;
			{8'd89, 8'd125}: color_data = 12'he01;
			{8'd89, 8'd126}: color_data = 12'he00;
			{8'd89, 8'd127}: color_data = 12'he00;
			{8'd89, 8'd128}: color_data = 12'he00;
			{8'd89, 8'd129}: color_data = 12'he00;
			{8'd89, 8'd130}: color_data = 12'he00;
			{8'd89, 8'd131}: color_data = 12'he00;
			{8'd89, 8'd132}: color_data = 12'he00;
			{8'd89, 8'd133}: color_data = 12'he00;
			{8'd89, 8'd134}: color_data = 12'hd00;
			{8'd89, 8'd138}: color_data = 12'he00;
			{8'd89, 8'd139}: color_data = 12'he00;
			{8'd89, 8'd140}: color_data = 12'he00;
			{8'd89, 8'd141}: color_data = 12'he00;
			{8'd89, 8'd142}: color_data = 12'he00;
			{8'd89, 8'd143}: color_data = 12'he01;
			{8'd89, 8'd144}: color_data = 12'he00;
			{8'd90, 8'd1}: color_data = 12'h000;
			{8'd90, 8'd2}: color_data = 12'h000;
			{8'd90, 8'd3}: color_data = 12'h000;
			{8'd90, 8'd4}: color_data = 12'h810;
			{8'd90, 8'd5}: color_data = 12'he21;
			{8'd90, 8'd6}: color_data = 12'he21;
			{8'd90, 8'd7}: color_data = 12'he21;
			{8'd90, 8'd8}: color_data = 12'he21;
			{8'd90, 8'd9}: color_data = 12'he21;
			{8'd90, 8'd10}: color_data = 12'he21;
			{8'd90, 8'd11}: color_data = 12'h710;
			{8'd90, 8'd12}: color_data = 12'h000;
			{8'd90, 8'd13}: color_data = 12'h000;
			{8'd90, 8'd14}: color_data = 12'h000;
			{8'd90, 8'd15}: color_data = 12'h000;
			{8'd90, 8'd16}: color_data = 12'h000;
			{8'd90, 8'd17}: color_data = 12'h200;
			{8'd90, 8'd18}: color_data = 12'he21;
			{8'd90, 8'd19}: color_data = 12'he21;
			{8'd90, 8'd20}: color_data = 12'he21;
			{8'd90, 8'd21}: color_data = 12'he21;
			{8'd90, 8'd22}: color_data = 12'he21;
			{8'd90, 8'd23}: color_data = 12'h810;
			{8'd90, 8'd24}: color_data = 12'h000;
			{8'd90, 8'd25}: color_data = 12'h000;
			{8'd90, 8'd26}: color_data = 12'h000;
			{8'd90, 8'd27}: color_data = 12'h000;
			{8'd90, 8'd28}: color_data = 12'h000;
			{8'd90, 8'd29}: color_data = 12'h000;
			{8'd90, 8'd30}: color_data = 12'h000;
			{8'd90, 8'd31}: color_data = 12'h000;
			{8'd90, 8'd32}: color_data = 12'h000;
			{8'd90, 8'd33}: color_data = 12'h000;
			{8'd90, 8'd34}: color_data = 12'heb0;
			{8'd90, 8'd35}: color_data = 12'hfd0;
			{8'd90, 8'd36}: color_data = 12'hfc0;
			{8'd90, 8'd37}: color_data = 12'hfc0;
			{8'd90, 8'd38}: color_data = 12'hfc0;
			{8'd90, 8'd39}: color_data = 12'hfc0;
			{8'd90, 8'd40}: color_data = 12'hfc0;
			{8'd90, 8'd41}: color_data = 12'hfd0;
			{8'd90, 8'd42}: color_data = 12'hfd0;
			{8'd90, 8'd43}: color_data = 12'hfd0;
			{8'd90, 8'd44}: color_data = 12'hfd0;
			{8'd90, 8'd45}: color_data = 12'hfd0;
			{8'd90, 8'd46}: color_data = 12'hfd0;
			{8'd90, 8'd47}: color_data = 12'hfd0;
			{8'd90, 8'd48}: color_data = 12'hfd0;
			{8'd90, 8'd49}: color_data = 12'hfd0;
			{8'd90, 8'd50}: color_data = 12'hfd0;
			{8'd90, 8'd51}: color_data = 12'hfd0;
			{8'd90, 8'd52}: color_data = 12'hfc0;
			{8'd90, 8'd53}: color_data = 12'hfc0;
			{8'd90, 8'd54}: color_data = 12'hfc0;
			{8'd90, 8'd55}: color_data = 12'hfc0;
			{8'd90, 8'd56}: color_data = 12'hfd0;
			{8'd90, 8'd57}: color_data = 12'hfd0;
			{8'd90, 8'd58}: color_data = 12'hfd0;
			{8'd90, 8'd59}: color_data = 12'hfd0;
			{8'd90, 8'd60}: color_data = 12'hfd0;
			{8'd90, 8'd61}: color_data = 12'hfd0;
			{8'd90, 8'd62}: color_data = 12'hfd0;
			{8'd90, 8'd63}: color_data = 12'hfd0;
			{8'd90, 8'd64}: color_data = 12'hfd0;
			{8'd90, 8'd65}: color_data = 12'hfd0;
			{8'd90, 8'd66}: color_data = 12'hfd0;
			{8'd90, 8'd67}: color_data = 12'h870;
			{8'd90, 8'd68}: color_data = 12'h000;
			{8'd90, 8'd69}: color_data = 12'h000;
			{8'd90, 8'd70}: color_data = 12'h000;
			{8'd90, 8'd71}: color_data = 12'h000;
			{8'd90, 8'd72}: color_data = 12'h000;
			{8'd90, 8'd73}: color_data = 12'h000;
			{8'd90, 8'd74}: color_data = 12'h000;
			{8'd90, 8'd100}: color_data = 12'he00;
			{8'd90, 8'd101}: color_data = 12'hf01;
			{8'd90, 8'd102}: color_data = 12'he00;
			{8'd90, 8'd103}: color_data = 12'he00;
			{8'd90, 8'd104}: color_data = 12'he00;
			{8'd90, 8'd105}: color_data = 12'he00;
			{8'd90, 8'd106}: color_data = 12'hc00;
			{8'd90, 8'd117}: color_data = 12'he00;
			{8'd90, 8'd118}: color_data = 12'he01;
			{8'd90, 8'd119}: color_data = 12'he00;
			{8'd90, 8'd120}: color_data = 12'he00;
			{8'd90, 8'd121}: color_data = 12'he00;
			{8'd90, 8'd124}: color_data = 12'he00;
			{8'd90, 8'd125}: color_data = 12'he00;
			{8'd90, 8'd126}: color_data = 12'he00;
			{8'd90, 8'd127}: color_data = 12'he00;
			{8'd90, 8'd130}: color_data = 12'he00;
			{8'd90, 8'd131}: color_data = 12'he01;
			{8'd90, 8'd132}: color_data = 12'he00;
			{8'd90, 8'd133}: color_data = 12'he00;
			{8'd90, 8'd138}: color_data = 12'he00;
			{8'd90, 8'd139}: color_data = 12'he00;
			{8'd90, 8'd140}: color_data = 12'he00;
			{8'd90, 8'd141}: color_data = 12'he00;
			{8'd90, 8'd142}: color_data = 12'he00;
			{8'd90, 8'd143}: color_data = 12'he01;
			{8'd90, 8'd144}: color_data = 12'he00;
			{8'd91, 8'd1}: color_data = 12'h000;
			{8'd91, 8'd2}: color_data = 12'h000;
			{8'd91, 8'd3}: color_data = 12'h000;
			{8'd91, 8'd4}: color_data = 12'h910;
			{8'd91, 8'd5}: color_data = 12'he21;
			{8'd91, 8'd6}: color_data = 12'he21;
			{8'd91, 8'd7}: color_data = 12'he21;
			{8'd91, 8'd8}: color_data = 12'he21;
			{8'd91, 8'd9}: color_data = 12'he21;
			{8'd91, 8'd10}: color_data = 12'he21;
			{8'd91, 8'd11}: color_data = 12'hc10;
			{8'd91, 8'd12}: color_data = 12'h000;
			{8'd91, 8'd13}: color_data = 12'h000;
			{8'd91, 8'd14}: color_data = 12'h000;
			{8'd91, 8'd15}: color_data = 12'h000;
			{8'd91, 8'd16}: color_data = 12'h000;
			{8'd91, 8'd17}: color_data = 12'h400;
			{8'd91, 8'd18}: color_data = 12'he21;
			{8'd91, 8'd19}: color_data = 12'he21;
			{8'd91, 8'd20}: color_data = 12'he21;
			{8'd91, 8'd21}: color_data = 12'he21;
			{8'd91, 8'd22}: color_data = 12'he21;
			{8'd91, 8'd23}: color_data = 12'h710;
			{8'd91, 8'd24}: color_data = 12'h000;
			{8'd91, 8'd25}: color_data = 12'h000;
			{8'd91, 8'd26}: color_data = 12'h000;
			{8'd91, 8'd27}: color_data = 12'h000;
			{8'd91, 8'd28}: color_data = 12'h000;
			{8'd91, 8'd29}: color_data = 12'h000;
			{8'd91, 8'd30}: color_data = 12'h000;
			{8'd91, 8'd31}: color_data = 12'h000;
			{8'd91, 8'd32}: color_data = 12'h000;
			{8'd91, 8'd33}: color_data = 12'h220;
			{8'd91, 8'd34}: color_data = 12'hfc0;
			{8'd91, 8'd35}: color_data = 12'hfd0;
			{8'd91, 8'd36}: color_data = 12'hfc0;
			{8'd91, 8'd37}: color_data = 12'hfc0;
			{8'd91, 8'd38}: color_data = 12'hfc0;
			{8'd91, 8'd39}: color_data = 12'hfc0;
			{8'd91, 8'd40}: color_data = 12'hfd0;
			{8'd91, 8'd41}: color_data = 12'hca0;
			{8'd91, 8'd42}: color_data = 12'h650;
			{8'd91, 8'd43}: color_data = 12'h750;
			{8'd91, 8'd44}: color_data = 12'h760;
			{8'd91, 8'd45}: color_data = 12'h860;
			{8'd91, 8'd46}: color_data = 12'h870;
			{8'd91, 8'd47}: color_data = 12'h970;
			{8'd91, 8'd48}: color_data = 12'h980;
			{8'd91, 8'd49}: color_data = 12'ha80;
			{8'd91, 8'd50}: color_data = 12'ha80;
			{8'd91, 8'd51}: color_data = 12'hdb0;
			{8'd91, 8'd52}: color_data = 12'hfd0;
			{8'd91, 8'd53}: color_data = 12'hfc0;
			{8'd91, 8'd54}: color_data = 12'hfc0;
			{8'd91, 8'd55}: color_data = 12'hfd0;
			{8'd91, 8'd56}: color_data = 12'heb0;
			{8'd91, 8'd57}: color_data = 12'hdb0;
			{8'd91, 8'd58}: color_data = 12'heb0;
			{8'd91, 8'd59}: color_data = 12'hec0;
			{8'd91, 8'd60}: color_data = 12'hec0;
			{8'd91, 8'd61}: color_data = 12'hfc0;
			{8'd91, 8'd62}: color_data = 12'hfc0;
			{8'd91, 8'd63}: color_data = 12'hfc0;
			{8'd91, 8'd64}: color_data = 12'hfd0;
			{8'd91, 8'd65}: color_data = 12'hfd0;
			{8'd91, 8'd66}: color_data = 12'hfd0;
			{8'd91, 8'd67}: color_data = 12'h760;
			{8'd91, 8'd68}: color_data = 12'h000;
			{8'd91, 8'd69}: color_data = 12'h000;
			{8'd91, 8'd70}: color_data = 12'h000;
			{8'd91, 8'd71}: color_data = 12'h000;
			{8'd91, 8'd72}: color_data = 12'h000;
			{8'd91, 8'd73}: color_data = 12'h000;
			{8'd91, 8'd74}: color_data = 12'h000;
			{8'd91, 8'd100}: color_data = 12'he00;
			{8'd91, 8'd101}: color_data = 12'hf01;
			{8'd91, 8'd102}: color_data = 12'he00;
			{8'd91, 8'd103}: color_data = 12'he00;
			{8'd91, 8'd104}: color_data = 12'he00;
			{8'd91, 8'd105}: color_data = 12'he00;
			{8'd91, 8'd106}: color_data = 12'hc00;
			{8'd91, 8'd117}: color_data = 12'he00;
			{8'd91, 8'd118}: color_data = 12'he01;
			{8'd91, 8'd119}: color_data = 12'he00;
			{8'd91, 8'd120}: color_data = 12'he00;
			{8'd91, 8'd121}: color_data = 12'he00;
			{8'd91, 8'd123}: color_data = 12'he00;
			{8'd91, 8'd124}: color_data = 12'he00;
			{8'd91, 8'd125}: color_data = 12'he00;
			{8'd91, 8'd126}: color_data = 12'he00;
			{8'd91, 8'd127}: color_data = 12'he00;
			{8'd91, 8'd130}: color_data = 12'he00;
			{8'd91, 8'd131}: color_data = 12'he01;
			{8'd91, 8'd132}: color_data = 12'he01;
			{8'd91, 8'd133}: color_data = 12'he00;
			{8'd91, 8'd138}: color_data = 12'he00;
			{8'd91, 8'd139}: color_data = 12'he00;
			{8'd91, 8'd140}: color_data = 12'he00;
			{8'd91, 8'd141}: color_data = 12'he00;
			{8'd91, 8'd142}: color_data = 12'he00;
			{8'd91, 8'd143}: color_data = 12'he01;
			{8'd91, 8'd144}: color_data = 12'he00;
			{8'd92, 8'd1}: color_data = 12'h000;
			{8'd92, 8'd2}: color_data = 12'h000;
			{8'd92, 8'd3}: color_data = 12'h000;
			{8'd92, 8'd4}: color_data = 12'h400;
			{8'd92, 8'd5}: color_data = 12'he21;
			{8'd92, 8'd6}: color_data = 12'he21;
			{8'd92, 8'd7}: color_data = 12'he21;
			{8'd92, 8'd8}: color_data = 12'he21;
			{8'd92, 8'd9}: color_data = 12'he21;
			{8'd92, 8'd10}: color_data = 12'he21;
			{8'd92, 8'd11}: color_data = 12'he21;
			{8'd92, 8'd12}: color_data = 12'h300;
			{8'd92, 8'd13}: color_data = 12'h000;
			{8'd92, 8'd14}: color_data = 12'h200;
			{8'd92, 8'd15}: color_data = 12'h400;
			{8'd92, 8'd16}: color_data = 12'h610;
			{8'd92, 8'd17}: color_data = 12'hb10;
			{8'd92, 8'd18}: color_data = 12'he21;
			{8'd92, 8'd19}: color_data = 12'he21;
			{8'd92, 8'd20}: color_data = 12'he21;
			{8'd92, 8'd21}: color_data = 12'he21;
			{8'd92, 8'd22}: color_data = 12'he21;
			{8'd92, 8'd23}: color_data = 12'h710;
			{8'd92, 8'd24}: color_data = 12'h000;
			{8'd92, 8'd25}: color_data = 12'h000;
			{8'd92, 8'd26}: color_data = 12'h000;
			{8'd92, 8'd27}: color_data = 12'h000;
			{8'd92, 8'd28}: color_data = 12'h000;
			{8'd92, 8'd29}: color_data = 12'h000;
			{8'd92, 8'd30}: color_data = 12'h000;
			{8'd92, 8'd31}: color_data = 12'h000;
			{8'd92, 8'd32}: color_data = 12'h000;
			{8'd92, 8'd33}: color_data = 12'h430;
			{8'd92, 8'd34}: color_data = 12'hfd0;
			{8'd92, 8'd35}: color_data = 12'hfc0;
			{8'd92, 8'd36}: color_data = 12'hfc0;
			{8'd92, 8'd37}: color_data = 12'hfc0;
			{8'd92, 8'd38}: color_data = 12'hfc0;
			{8'd92, 8'd39}: color_data = 12'hfc0;
			{8'd92, 8'd40}: color_data = 12'hfd0;
			{8'd92, 8'd41}: color_data = 12'hda0;
			{8'd92, 8'd42}: color_data = 12'h000;
			{8'd92, 8'd43}: color_data = 12'h000;
			{8'd92, 8'd44}: color_data = 12'h000;
			{8'd92, 8'd45}: color_data = 12'h000;
			{8'd92, 8'd46}: color_data = 12'h000;
			{8'd92, 8'd47}: color_data = 12'h000;
			{8'd92, 8'd48}: color_data = 12'h000;
			{8'd92, 8'd49}: color_data = 12'h000;
			{8'd92, 8'd50}: color_data = 12'h000;
			{8'd92, 8'd51}: color_data = 12'hb90;
			{8'd92, 8'd52}: color_data = 12'hfd0;
			{8'd92, 8'd53}: color_data = 12'hfc0;
			{8'd92, 8'd54}: color_data = 12'hfc0;
			{8'd92, 8'd55}: color_data = 12'hfd0;
			{8'd92, 8'd56}: color_data = 12'hca0;
			{8'd92, 8'd57}: color_data = 12'h220;
			{8'd92, 8'd58}: color_data = 12'h000;
			{8'd92, 8'd59}: color_data = 12'h110;
			{8'd92, 8'd60}: color_data = 12'h110;
			{8'd92, 8'd61}: color_data = 12'h210;
			{8'd92, 8'd62}: color_data = 12'h220;
			{8'd92, 8'd63}: color_data = 12'h320;
			{8'd92, 8'd64}: color_data = 12'h320;
			{8'd92, 8'd65}: color_data = 12'h430;
			{8'd92, 8'd66}: color_data = 12'h430;
			{8'd92, 8'd67}: color_data = 12'h110;
			{8'd92, 8'd68}: color_data = 12'h000;
			{8'd92, 8'd69}: color_data = 12'h000;
			{8'd92, 8'd70}: color_data = 12'h000;
			{8'd92, 8'd71}: color_data = 12'h000;
			{8'd92, 8'd72}: color_data = 12'h000;
			{8'd92, 8'd73}: color_data = 12'h000;
			{8'd92, 8'd74}: color_data = 12'h000;
			{8'd92, 8'd100}: color_data = 12'he00;
			{8'd92, 8'd101}: color_data = 12'hf01;
			{8'd92, 8'd102}: color_data = 12'he00;
			{8'd92, 8'd103}: color_data = 12'he00;
			{8'd92, 8'd104}: color_data = 12'he00;
			{8'd92, 8'd105}: color_data = 12'he00;
			{8'd92, 8'd106}: color_data = 12'hc00;
			{8'd92, 8'd117}: color_data = 12'he00;
			{8'd92, 8'd118}: color_data = 12'he01;
			{8'd92, 8'd119}: color_data = 12'he00;
			{8'd92, 8'd120}: color_data = 12'he00;
			{8'd92, 8'd121}: color_data = 12'he00;
			{8'd92, 8'd123}: color_data = 12'he01;
			{8'd92, 8'd124}: color_data = 12'he00;
			{8'd92, 8'd125}: color_data = 12'he01;
			{8'd92, 8'd126}: color_data = 12'he00;
			{8'd92, 8'd130}: color_data = 12'he00;
			{8'd92, 8'd131}: color_data = 12'he01;
			{8'd92, 8'd132}: color_data = 12'he00;
			{8'd92, 8'd133}: color_data = 12'he00;
			{8'd92, 8'd138}: color_data = 12'he00;
			{8'd92, 8'd139}: color_data = 12'he00;
			{8'd92, 8'd140}: color_data = 12'he00;
			{8'd92, 8'd141}: color_data = 12'he00;
			{8'd92, 8'd142}: color_data = 12'he00;
			{8'd92, 8'd143}: color_data = 12'he01;
			{8'd92, 8'd144}: color_data = 12'he00;
			{8'd93, 8'd2}: color_data = 12'h000;
			{8'd93, 8'd3}: color_data = 12'h000;
			{8'd93, 8'd4}: color_data = 12'h000;
			{8'd93, 8'd5}: color_data = 12'ha10;
			{8'd93, 8'd6}: color_data = 12'he21;
			{8'd93, 8'd7}: color_data = 12'he21;
			{8'd93, 8'd8}: color_data = 12'he21;
			{8'd93, 8'd9}: color_data = 12'he21;
			{8'd93, 8'd10}: color_data = 12'he21;
			{8'd93, 8'd11}: color_data = 12'he21;
			{8'd93, 8'd12}: color_data = 12'hd20;
			{8'd93, 8'd13}: color_data = 12'hd20;
			{8'd93, 8'd14}: color_data = 12'he21;
			{8'd93, 8'd15}: color_data = 12'he21;
			{8'd93, 8'd16}: color_data = 12'hf21;
			{8'd93, 8'd17}: color_data = 12'he21;
			{8'd93, 8'd18}: color_data = 12'he21;
			{8'd93, 8'd19}: color_data = 12'he21;
			{8'd93, 8'd20}: color_data = 12'he21;
			{8'd93, 8'd21}: color_data = 12'he21;
			{8'd93, 8'd22}: color_data = 12'hf21;
			{8'd93, 8'd23}: color_data = 12'h600;
			{8'd93, 8'd24}: color_data = 12'h000;
			{8'd93, 8'd25}: color_data = 12'h000;
			{8'd93, 8'd26}: color_data = 12'h000;
			{8'd93, 8'd27}: color_data = 12'h000;
			{8'd93, 8'd28}: color_data = 12'h000;
			{8'd93, 8'd29}: color_data = 12'h000;
			{8'd93, 8'd30}: color_data = 12'h000;
			{8'd93, 8'd31}: color_data = 12'h000;
			{8'd93, 8'd32}: color_data = 12'h000;
			{8'd93, 8'd33}: color_data = 12'h650;
			{8'd93, 8'd34}: color_data = 12'hfd0;
			{8'd93, 8'd35}: color_data = 12'hfc0;
			{8'd93, 8'd36}: color_data = 12'hfc0;
			{8'd93, 8'd37}: color_data = 12'hfc0;
			{8'd93, 8'd38}: color_data = 12'hfc0;
			{8'd93, 8'd39}: color_data = 12'hfc0;
			{8'd93, 8'd40}: color_data = 12'hfd0;
			{8'd93, 8'd41}: color_data = 12'hfc0;
			{8'd93, 8'd42}: color_data = 12'h320;
			{8'd93, 8'd43}: color_data = 12'h000;
			{8'd93, 8'd44}: color_data = 12'h000;
			{8'd93, 8'd45}: color_data = 12'h000;
			{8'd93, 8'd46}: color_data = 12'h000;
			{8'd93, 8'd47}: color_data = 12'h000;
			{8'd93, 8'd48}: color_data = 12'h000;
			{8'd93, 8'd49}: color_data = 12'h000;
			{8'd93, 8'd50}: color_data = 12'h100;
			{8'd93, 8'd51}: color_data = 12'hdb0;
			{8'd93, 8'd52}: color_data = 12'hfd0;
			{8'd93, 8'd53}: color_data = 12'hfc0;
			{8'd93, 8'd54}: color_data = 12'hfc0;
			{8'd93, 8'd55}: color_data = 12'hfc0;
			{8'd93, 8'd56}: color_data = 12'hfd0;
			{8'd93, 8'd57}: color_data = 12'heb0;
			{8'd93, 8'd58}: color_data = 12'h540;
			{8'd93, 8'd59}: color_data = 12'h000;
			{8'd93, 8'd60}: color_data = 12'h000;
			{8'd93, 8'd61}: color_data = 12'h000;
			{8'd93, 8'd62}: color_data = 12'h000;
			{8'd93, 8'd63}: color_data = 12'h000;
			{8'd93, 8'd64}: color_data = 12'h000;
			{8'd93, 8'd65}: color_data = 12'h000;
			{8'd93, 8'd66}: color_data = 12'h000;
			{8'd93, 8'd67}: color_data = 12'h000;
			{8'd93, 8'd68}: color_data = 12'h000;
			{8'd93, 8'd69}: color_data = 12'h000;
			{8'd93, 8'd70}: color_data = 12'h000;
			{8'd93, 8'd71}: color_data = 12'h000;
			{8'd93, 8'd72}: color_data = 12'h000;
			{8'd93, 8'd73}: color_data = 12'h000;
			{8'd93, 8'd74}: color_data = 12'h000;
			{8'd93, 8'd100}: color_data = 12'he00;
			{8'd93, 8'd101}: color_data = 12'hf01;
			{8'd93, 8'd102}: color_data = 12'he00;
			{8'd93, 8'd103}: color_data = 12'he00;
			{8'd93, 8'd104}: color_data = 12'he00;
			{8'd93, 8'd105}: color_data = 12'he00;
			{8'd93, 8'd106}: color_data = 12'hc00;
			{8'd93, 8'd117}: color_data = 12'he00;
			{8'd93, 8'd118}: color_data = 12'he01;
			{8'd93, 8'd119}: color_data = 12'he00;
			{8'd93, 8'd120}: color_data = 12'he00;
			{8'd93, 8'd121}: color_data = 12'he00;
			{8'd93, 8'd123}: color_data = 12'he00;
			{8'd93, 8'd124}: color_data = 12'he01;
			{8'd93, 8'd125}: color_data = 12'he01;
			{8'd93, 8'd126}: color_data = 12'he00;
			{8'd93, 8'd129}: color_data = 12'he00;
			{8'd93, 8'd130}: color_data = 12'he00;
			{8'd93, 8'd131}: color_data = 12'he01;
			{8'd93, 8'd132}: color_data = 12'he00;
			{8'd93, 8'd133}: color_data = 12'hf00;
			{8'd93, 8'd138}: color_data = 12'he00;
			{8'd93, 8'd139}: color_data = 12'he00;
			{8'd93, 8'd140}: color_data = 12'he00;
			{8'd93, 8'd141}: color_data = 12'he00;
			{8'd93, 8'd142}: color_data = 12'he00;
			{8'd93, 8'd143}: color_data = 12'he01;
			{8'd93, 8'd144}: color_data = 12'he00;
			{8'd94, 8'd2}: color_data = 12'h000;
			{8'd94, 8'd3}: color_data = 12'h000;
			{8'd94, 8'd4}: color_data = 12'h000;
			{8'd94, 8'd5}: color_data = 12'h300;
			{8'd94, 8'd6}: color_data = 12'he21;
			{8'd94, 8'd7}: color_data = 12'he21;
			{8'd94, 8'd8}: color_data = 12'he21;
			{8'd94, 8'd9}: color_data = 12'he21;
			{8'd94, 8'd10}: color_data = 12'he21;
			{8'd94, 8'd11}: color_data = 12'he21;
			{8'd94, 8'd12}: color_data = 12'he21;
			{8'd94, 8'd13}: color_data = 12'he21;
			{8'd94, 8'd14}: color_data = 12'he21;
			{8'd94, 8'd15}: color_data = 12'he21;
			{8'd94, 8'd16}: color_data = 12'he21;
			{8'd94, 8'd17}: color_data = 12'he21;
			{8'd94, 8'd18}: color_data = 12'he21;
			{8'd94, 8'd19}: color_data = 12'he21;
			{8'd94, 8'd20}: color_data = 12'he21;
			{8'd94, 8'd21}: color_data = 12'he21;
			{8'd94, 8'd22}: color_data = 12'hd21;
			{8'd94, 8'd23}: color_data = 12'h200;
			{8'd94, 8'd24}: color_data = 12'h000;
			{8'd94, 8'd25}: color_data = 12'h000;
			{8'd94, 8'd26}: color_data = 12'h000;
			{8'd94, 8'd27}: color_data = 12'h000;
			{8'd94, 8'd28}: color_data = 12'h000;
			{8'd94, 8'd29}: color_data = 12'h000;
			{8'd94, 8'd30}: color_data = 12'h000;
			{8'd94, 8'd31}: color_data = 12'h000;
			{8'd94, 8'd32}: color_data = 12'h000;
			{8'd94, 8'd33}: color_data = 12'h970;
			{8'd94, 8'd34}: color_data = 12'hfd0;
			{8'd94, 8'd35}: color_data = 12'hfc0;
			{8'd94, 8'd36}: color_data = 12'hfc0;
			{8'd94, 8'd37}: color_data = 12'hfc0;
			{8'd94, 8'd38}: color_data = 12'hfc0;
			{8'd94, 8'd39}: color_data = 12'hfc0;
			{8'd94, 8'd40}: color_data = 12'hfc0;
			{8'd94, 8'd41}: color_data = 12'hfd0;
			{8'd94, 8'd42}: color_data = 12'h650;
			{8'd94, 8'd43}: color_data = 12'h000;
			{8'd94, 8'd44}: color_data = 12'h000;
			{8'd94, 8'd45}: color_data = 12'h000;
			{8'd94, 8'd46}: color_data = 12'h000;
			{8'd94, 8'd47}: color_data = 12'h000;
			{8'd94, 8'd48}: color_data = 12'h000;
			{8'd94, 8'd49}: color_data = 12'h000;
			{8'd94, 8'd50}: color_data = 12'h320;
			{8'd94, 8'd51}: color_data = 12'hfc0;
			{8'd94, 8'd52}: color_data = 12'hfd0;
			{8'd94, 8'd53}: color_data = 12'hfc0;
			{8'd94, 8'd54}: color_data = 12'hfc0;
			{8'd94, 8'd55}: color_data = 12'hfc0;
			{8'd94, 8'd56}: color_data = 12'hfc0;
			{8'd94, 8'd57}: color_data = 12'hfd0;
			{8'd94, 8'd58}: color_data = 12'hfd0;
			{8'd94, 8'd59}: color_data = 12'ha80;
			{8'd94, 8'd60}: color_data = 12'h210;
			{8'd94, 8'd61}: color_data = 12'h000;
			{8'd94, 8'd62}: color_data = 12'h000;
			{8'd94, 8'd63}: color_data = 12'h000;
			{8'd94, 8'd64}: color_data = 12'h000;
			{8'd94, 8'd65}: color_data = 12'h000;
			{8'd94, 8'd66}: color_data = 12'h000;
			{8'd94, 8'd67}: color_data = 12'h000;
			{8'd94, 8'd68}: color_data = 12'h000;
			{8'd94, 8'd69}: color_data = 12'h000;
			{8'd94, 8'd70}: color_data = 12'h000;
			{8'd94, 8'd71}: color_data = 12'h000;
			{8'd94, 8'd72}: color_data = 12'h000;
			{8'd94, 8'd73}: color_data = 12'h000;
			{8'd94, 8'd74}: color_data = 12'h000;
			{8'd94, 8'd100}: color_data = 12'he00;
			{8'd94, 8'd101}: color_data = 12'hf01;
			{8'd94, 8'd102}: color_data = 12'he00;
			{8'd94, 8'd103}: color_data = 12'he00;
			{8'd94, 8'd104}: color_data = 12'he00;
			{8'd94, 8'd105}: color_data = 12'he00;
			{8'd94, 8'd106}: color_data = 12'hc00;
			{8'd94, 8'd117}: color_data = 12'he00;
			{8'd94, 8'd118}: color_data = 12'he01;
			{8'd94, 8'd119}: color_data = 12'he00;
			{8'd94, 8'd120}: color_data = 12'he00;
			{8'd94, 8'd121}: color_data = 12'he00;
			{8'd94, 8'd122}: color_data = 12'he00;
			{8'd94, 8'd123}: color_data = 12'he00;
			{8'd94, 8'd124}: color_data = 12'he00;
			{8'd94, 8'd125}: color_data = 12'he00;
			{8'd94, 8'd126}: color_data = 12'he00;
			{8'd94, 8'd127}: color_data = 12'he01;
			{8'd94, 8'd128}: color_data = 12'he00;
			{8'd94, 8'd129}: color_data = 12'he00;
			{8'd94, 8'd130}: color_data = 12'he00;
			{8'd94, 8'd131}: color_data = 12'he00;
			{8'd94, 8'd132}: color_data = 12'he00;
			{8'd94, 8'd138}: color_data = 12'he00;
			{8'd94, 8'd139}: color_data = 12'he00;
			{8'd94, 8'd140}: color_data = 12'he00;
			{8'd94, 8'd141}: color_data = 12'he00;
			{8'd94, 8'd142}: color_data = 12'he00;
			{8'd94, 8'd143}: color_data = 12'he01;
			{8'd94, 8'd144}: color_data = 12'he00;
			{8'd95, 8'd3}: color_data = 12'h000;
			{8'd95, 8'd4}: color_data = 12'h000;
			{8'd95, 8'd5}: color_data = 12'h000;
			{8'd95, 8'd6}: color_data = 12'h910;
			{8'd95, 8'd7}: color_data = 12'he21;
			{8'd95, 8'd8}: color_data = 12'he21;
			{8'd95, 8'd9}: color_data = 12'he21;
			{8'd95, 8'd10}: color_data = 12'he21;
			{8'd95, 8'd11}: color_data = 12'he21;
			{8'd95, 8'd12}: color_data = 12'he21;
			{8'd95, 8'd13}: color_data = 12'he21;
			{8'd95, 8'd14}: color_data = 12'he21;
			{8'd95, 8'd15}: color_data = 12'he21;
			{8'd95, 8'd16}: color_data = 12'he21;
			{8'd95, 8'd17}: color_data = 12'he21;
			{8'd95, 8'd18}: color_data = 12'he21;
			{8'd95, 8'd19}: color_data = 12'he21;
			{8'd95, 8'd20}: color_data = 12'he21;
			{8'd95, 8'd21}: color_data = 12'he20;
			{8'd95, 8'd22}: color_data = 12'h400;
			{8'd95, 8'd23}: color_data = 12'h000;
			{8'd95, 8'd24}: color_data = 12'h000;
			{8'd95, 8'd25}: color_data = 12'h000;
			{8'd95, 8'd26}: color_data = 12'h000;
			{8'd95, 8'd27}: color_data = 12'h000;
			{8'd95, 8'd28}: color_data = 12'h000;
			{8'd95, 8'd29}: color_data = 12'h000;
			{8'd95, 8'd30}: color_data = 12'h000;
			{8'd95, 8'd31}: color_data = 12'h000;
			{8'd95, 8'd32}: color_data = 12'h000;
			{8'd95, 8'd33}: color_data = 12'hb90;
			{8'd95, 8'd34}: color_data = 12'hfd0;
			{8'd95, 8'd35}: color_data = 12'hfc0;
			{8'd95, 8'd36}: color_data = 12'hfc0;
			{8'd95, 8'd37}: color_data = 12'hfc0;
			{8'd95, 8'd38}: color_data = 12'hfc0;
			{8'd95, 8'd39}: color_data = 12'hfc0;
			{8'd95, 8'd40}: color_data = 12'hfc0;
			{8'd95, 8'd41}: color_data = 12'hfd0;
			{8'd95, 8'd42}: color_data = 12'hb90;
			{8'd95, 8'd43}: color_data = 12'h000;
			{8'd95, 8'd44}: color_data = 12'h000;
			{8'd95, 8'd45}: color_data = 12'h000;
			{8'd95, 8'd46}: color_data = 12'h000;
			{8'd95, 8'd47}: color_data = 12'h000;
			{8'd95, 8'd48}: color_data = 12'h000;
			{8'd95, 8'd49}: color_data = 12'h000;
			{8'd95, 8'd50}: color_data = 12'h650;
			{8'd95, 8'd51}: color_data = 12'hfd0;
			{8'd95, 8'd52}: color_data = 12'hfc0;
			{8'd95, 8'd53}: color_data = 12'hfc0;
			{8'd95, 8'd54}: color_data = 12'hfc0;
			{8'd95, 8'd55}: color_data = 12'hfc0;
			{8'd95, 8'd56}: color_data = 12'hfc0;
			{8'd95, 8'd57}: color_data = 12'hfc0;
			{8'd95, 8'd58}: color_data = 12'hfd0;
			{8'd95, 8'd59}: color_data = 12'hfd0;
			{8'd95, 8'd60}: color_data = 12'heb0;
			{8'd95, 8'd61}: color_data = 12'h650;
			{8'd95, 8'd62}: color_data = 12'h000;
			{8'd95, 8'd63}: color_data = 12'h000;
			{8'd95, 8'd64}: color_data = 12'h000;
			{8'd95, 8'd65}: color_data = 12'h000;
			{8'd95, 8'd66}: color_data = 12'h000;
			{8'd95, 8'd67}: color_data = 12'h000;
			{8'd95, 8'd68}: color_data = 12'h000;
			{8'd95, 8'd69}: color_data = 12'h000;
			{8'd95, 8'd70}: color_data = 12'h000;
			{8'd95, 8'd71}: color_data = 12'h000;
			{8'd95, 8'd72}: color_data = 12'h000;
			{8'd95, 8'd73}: color_data = 12'h000;
			{8'd95, 8'd100}: color_data = 12'he00;
			{8'd95, 8'd101}: color_data = 12'hf01;
			{8'd95, 8'd102}: color_data = 12'he00;
			{8'd95, 8'd103}: color_data = 12'he00;
			{8'd95, 8'd104}: color_data = 12'he00;
			{8'd95, 8'd105}: color_data = 12'he00;
			{8'd95, 8'd106}: color_data = 12'hc00;
			{8'd95, 8'd117}: color_data = 12'he00;
			{8'd95, 8'd118}: color_data = 12'he00;
			{8'd95, 8'd119}: color_data = 12'he00;
			{8'd95, 8'd120}: color_data = 12'he00;
			{8'd95, 8'd121}: color_data = 12'he01;
			{8'd95, 8'd122}: color_data = 12'he00;
			{8'd95, 8'd123}: color_data = 12'he00;
			{8'd95, 8'd124}: color_data = 12'he00;
			{8'd95, 8'd125}: color_data = 12'he00;
			{8'd95, 8'd126}: color_data = 12'he00;
			{8'd95, 8'd127}: color_data = 12'he00;
			{8'd95, 8'd128}: color_data = 12'he01;
			{8'd95, 8'd129}: color_data = 12'he00;
			{8'd95, 8'd130}: color_data = 12'he00;
			{8'd95, 8'd131}: color_data = 12'he00;
			{8'd95, 8'd132}: color_data = 12'he00;
			{8'd95, 8'd133}: color_data = 12'he00;
			{8'd95, 8'd138}: color_data = 12'he00;
			{8'd95, 8'd139}: color_data = 12'he00;
			{8'd95, 8'd140}: color_data = 12'he00;
			{8'd95, 8'd141}: color_data = 12'he00;
			{8'd95, 8'd142}: color_data = 12'he00;
			{8'd95, 8'd143}: color_data = 12'he01;
			{8'd95, 8'd144}: color_data = 12'he00;
			{8'd96, 8'd4}: color_data = 12'h000;
			{8'd96, 8'd5}: color_data = 12'h000;
			{8'd96, 8'd6}: color_data = 12'h200;
			{8'd96, 8'd7}: color_data = 12'hd20;
			{8'd96, 8'd8}: color_data = 12'he21;
			{8'd96, 8'd9}: color_data = 12'he21;
			{8'd96, 8'd10}: color_data = 12'he21;
			{8'd96, 8'd11}: color_data = 12'he21;
			{8'd96, 8'd12}: color_data = 12'he21;
			{8'd96, 8'd13}: color_data = 12'he21;
			{8'd96, 8'd14}: color_data = 12'he21;
			{8'd96, 8'd15}: color_data = 12'he21;
			{8'd96, 8'd16}: color_data = 12'he21;
			{8'd96, 8'd17}: color_data = 12'he21;
			{8'd96, 8'd18}: color_data = 12'he21;
			{8'd96, 8'd19}: color_data = 12'he21;
			{8'd96, 8'd20}: color_data = 12'he21;
			{8'd96, 8'd21}: color_data = 12'h400;
			{8'd96, 8'd22}: color_data = 12'h000;
			{8'd96, 8'd23}: color_data = 12'h000;
			{8'd96, 8'd24}: color_data = 12'h000;
			{8'd96, 8'd25}: color_data = 12'h000;
			{8'd96, 8'd26}: color_data = 12'h000;
			{8'd96, 8'd27}: color_data = 12'h000;
			{8'd96, 8'd28}: color_data = 12'h000;
			{8'd96, 8'd29}: color_data = 12'h000;
			{8'd96, 8'd30}: color_data = 12'h000;
			{8'd96, 8'd31}: color_data = 12'h000;
			{8'd96, 8'd32}: color_data = 12'h000;
			{8'd96, 8'd33}: color_data = 12'hdb0;
			{8'd96, 8'd34}: color_data = 12'hfd0;
			{8'd96, 8'd35}: color_data = 12'hfc0;
			{8'd96, 8'd36}: color_data = 12'hfc0;
			{8'd96, 8'd37}: color_data = 12'hfc0;
			{8'd96, 8'd38}: color_data = 12'hfc0;
			{8'd96, 8'd39}: color_data = 12'hfc0;
			{8'd96, 8'd40}: color_data = 12'hfc0;
			{8'd96, 8'd41}: color_data = 12'hfd0;
			{8'd96, 8'd42}: color_data = 12'heb0;
			{8'd96, 8'd43}: color_data = 12'h110;
			{8'd96, 8'd44}: color_data = 12'h000;
			{8'd96, 8'd45}: color_data = 12'h000;
			{8'd96, 8'd46}: color_data = 12'h000;
			{8'd96, 8'd47}: color_data = 12'h000;
			{8'd96, 8'd48}: color_data = 12'h000;
			{8'd96, 8'd49}: color_data = 12'h000;
			{8'd96, 8'd50}: color_data = 12'ha80;
			{8'd96, 8'd51}: color_data = 12'hfd0;
			{8'd96, 8'd52}: color_data = 12'hfc0;
			{8'd96, 8'd53}: color_data = 12'hfc0;
			{8'd96, 8'd54}: color_data = 12'hfc0;
			{8'd96, 8'd55}: color_data = 12'hfc0;
			{8'd96, 8'd56}: color_data = 12'hfc0;
			{8'd96, 8'd57}: color_data = 12'hfc0;
			{8'd96, 8'd58}: color_data = 12'hfc0;
			{8'd96, 8'd59}: color_data = 12'hfc0;
			{8'd96, 8'd60}: color_data = 12'hfd0;
			{8'd96, 8'd61}: color_data = 12'hfd0;
			{8'd96, 8'd62}: color_data = 12'hb90;
			{8'd96, 8'd63}: color_data = 12'h220;
			{8'd96, 8'd64}: color_data = 12'h000;
			{8'd96, 8'd65}: color_data = 12'h000;
			{8'd96, 8'd66}: color_data = 12'h000;
			{8'd96, 8'd67}: color_data = 12'h000;
			{8'd96, 8'd68}: color_data = 12'h000;
			{8'd96, 8'd69}: color_data = 12'h000;
			{8'd96, 8'd70}: color_data = 12'h000;
			{8'd96, 8'd71}: color_data = 12'h000;
			{8'd96, 8'd72}: color_data = 12'h000;
			{8'd96, 8'd100}: color_data = 12'he00;
			{8'd96, 8'd101}: color_data = 12'hf01;
			{8'd96, 8'd102}: color_data = 12'he00;
			{8'd96, 8'd103}: color_data = 12'he00;
			{8'd96, 8'd104}: color_data = 12'he00;
			{8'd96, 8'd105}: color_data = 12'he00;
			{8'd96, 8'd106}: color_data = 12'hc00;
			{8'd96, 8'd117}: color_data = 12'he01;
			{8'd96, 8'd118}: color_data = 12'he00;
			{8'd96, 8'd119}: color_data = 12'he00;
			{8'd96, 8'd120}: color_data = 12'he00;
			{8'd96, 8'd121}: color_data = 12'he00;
			{8'd96, 8'd122}: color_data = 12'he00;
			{8'd96, 8'd123}: color_data = 12'he00;
			{8'd96, 8'd124}: color_data = 12'he00;
			{8'd96, 8'd125}: color_data = 12'he00;
			{8'd96, 8'd126}: color_data = 12'he00;
			{8'd96, 8'd127}: color_data = 12'he00;
			{8'd96, 8'd128}: color_data = 12'he00;
			{8'd96, 8'd129}: color_data = 12'he00;
			{8'd96, 8'd130}: color_data = 12'he00;
			{8'd96, 8'd131}: color_data = 12'he00;
			{8'd96, 8'd132}: color_data = 12'hf01;
			{8'd96, 8'd133}: color_data = 12'he00;
			{8'd96, 8'd138}: color_data = 12'he00;
			{8'd96, 8'd139}: color_data = 12'he00;
			{8'd96, 8'd140}: color_data = 12'he00;
			{8'd96, 8'd141}: color_data = 12'he00;
			{8'd96, 8'd142}: color_data = 12'he00;
			{8'd96, 8'd143}: color_data = 12'he01;
			{8'd96, 8'd144}: color_data = 12'he00;
			{8'd97, 8'd4}: color_data = 12'h000;
			{8'd97, 8'd5}: color_data = 12'h000;
			{8'd97, 8'd6}: color_data = 12'h000;
			{8'd97, 8'd7}: color_data = 12'h810;
			{8'd97, 8'd8}: color_data = 12'hf21;
			{8'd97, 8'd9}: color_data = 12'he21;
			{8'd97, 8'd10}: color_data = 12'he21;
			{8'd97, 8'd11}: color_data = 12'he21;
			{8'd97, 8'd12}: color_data = 12'he21;
			{8'd97, 8'd13}: color_data = 12'he21;
			{8'd97, 8'd14}: color_data = 12'he21;
			{8'd97, 8'd15}: color_data = 12'he21;
			{8'd97, 8'd16}: color_data = 12'he21;
			{8'd97, 8'd17}: color_data = 12'he21;
			{8'd97, 8'd18}: color_data = 12'he21;
			{8'd97, 8'd19}: color_data = 12'he21;
			{8'd97, 8'd20}: color_data = 12'h500;
			{8'd97, 8'd21}: color_data = 12'h000;
			{8'd97, 8'd22}: color_data = 12'h000;
			{8'd97, 8'd23}: color_data = 12'h000;
			{8'd97, 8'd24}: color_data = 12'h000;
			{8'd97, 8'd25}: color_data = 12'h000;
			{8'd97, 8'd26}: color_data = 12'h000;
			{8'd97, 8'd27}: color_data = 12'h000;
			{8'd97, 8'd28}: color_data = 12'h000;
			{8'd97, 8'd29}: color_data = 12'h000;
			{8'd97, 8'd30}: color_data = 12'h000;
			{8'd97, 8'd31}: color_data = 12'h000;
			{8'd97, 8'd32}: color_data = 12'h000;
			{8'd97, 8'd33}: color_data = 12'hca0;
			{8'd97, 8'd34}: color_data = 12'hfd0;
			{8'd97, 8'd35}: color_data = 12'hfc0;
			{8'd97, 8'd36}: color_data = 12'hfc0;
			{8'd97, 8'd37}: color_data = 12'hfc0;
			{8'd97, 8'd38}: color_data = 12'hfc0;
			{8'd97, 8'd39}: color_data = 12'hfc0;
			{8'd97, 8'd40}: color_data = 12'hfc0;
			{8'd97, 8'd41}: color_data = 12'hfd0;
			{8'd97, 8'd42}: color_data = 12'hfd0;
			{8'd97, 8'd43}: color_data = 12'h430;
			{8'd97, 8'd44}: color_data = 12'h000;
			{8'd97, 8'd45}: color_data = 12'h000;
			{8'd97, 8'd46}: color_data = 12'h000;
			{8'd97, 8'd47}: color_data = 12'h000;
			{8'd97, 8'd48}: color_data = 12'h000;
			{8'd97, 8'd49}: color_data = 12'h220;
			{8'd97, 8'd50}: color_data = 12'hdb0;
			{8'd97, 8'd51}: color_data = 12'hfd0;
			{8'd97, 8'd52}: color_data = 12'hfc0;
			{8'd97, 8'd53}: color_data = 12'hfc0;
			{8'd97, 8'd54}: color_data = 12'hfc0;
			{8'd97, 8'd55}: color_data = 12'hfc0;
			{8'd97, 8'd56}: color_data = 12'hfc0;
			{8'd97, 8'd57}: color_data = 12'hfc0;
			{8'd97, 8'd58}: color_data = 12'hfc0;
			{8'd97, 8'd59}: color_data = 12'hfc0;
			{8'd97, 8'd60}: color_data = 12'hfc0;
			{8'd97, 8'd61}: color_data = 12'hfc0;
			{8'd97, 8'd62}: color_data = 12'hfd0;
			{8'd97, 8'd63}: color_data = 12'hec0;
			{8'd97, 8'd64}: color_data = 12'h650;
			{8'd97, 8'd65}: color_data = 12'h000;
			{8'd97, 8'd66}: color_data = 12'h000;
			{8'd97, 8'd67}: color_data = 12'h000;
			{8'd97, 8'd68}: color_data = 12'h000;
			{8'd97, 8'd69}: color_data = 12'h000;
			{8'd97, 8'd70}: color_data = 12'h000;
			{8'd97, 8'd71}: color_data = 12'h000;
			{8'd97, 8'd72}: color_data = 12'h000;
			{8'd97, 8'd73}: color_data = 12'h000;
			{8'd97, 8'd74}: color_data = 12'h000;
			{8'd97, 8'd100}: color_data = 12'he00;
			{8'd97, 8'd101}: color_data = 12'hf01;
			{8'd97, 8'd102}: color_data = 12'he00;
			{8'd97, 8'd103}: color_data = 12'he00;
			{8'd97, 8'd104}: color_data = 12'he00;
			{8'd97, 8'd105}: color_data = 12'he00;
			{8'd97, 8'd106}: color_data = 12'hc00;
			{8'd97, 8'd117}: color_data = 12'ha00;
			{8'd97, 8'd118}: color_data = 12'he00;
			{8'd97, 8'd119}: color_data = 12'he00;
			{8'd97, 8'd120}: color_data = 12'he00;
			{8'd97, 8'd121}: color_data = 12'he00;
			{8'd97, 8'd122}: color_data = 12'he00;
			{8'd97, 8'd123}: color_data = 12'he00;
			{8'd97, 8'd124}: color_data = 12'he00;
			{8'd97, 8'd125}: color_data = 12'he00;
			{8'd97, 8'd126}: color_data = 12'he00;
			{8'd97, 8'd127}: color_data = 12'he00;
			{8'd97, 8'd128}: color_data = 12'he00;
			{8'd97, 8'd129}: color_data = 12'he00;
			{8'd97, 8'd130}: color_data = 12'he00;
			{8'd97, 8'd131}: color_data = 12'he00;
			{8'd97, 8'd132}: color_data = 12'hf01;
			{8'd97, 8'd133}: color_data = 12'he00;
			{8'd97, 8'd138}: color_data = 12'he00;
			{8'd97, 8'd139}: color_data = 12'he00;
			{8'd97, 8'd140}: color_data = 12'he00;
			{8'd97, 8'd141}: color_data = 12'he00;
			{8'd97, 8'd142}: color_data = 12'he00;
			{8'd97, 8'd143}: color_data = 12'he01;
			{8'd97, 8'd144}: color_data = 12'he00;
			{8'd98, 8'd5}: color_data = 12'h000;
			{8'd98, 8'd6}: color_data = 12'h000;
			{8'd98, 8'd7}: color_data = 12'h100;
			{8'd98, 8'd8}: color_data = 12'hd20;
			{8'd98, 8'd9}: color_data = 12'he21;
			{8'd98, 8'd10}: color_data = 12'he21;
			{8'd98, 8'd11}: color_data = 12'he21;
			{8'd98, 8'd12}: color_data = 12'he21;
			{8'd98, 8'd13}: color_data = 12'he21;
			{8'd98, 8'd14}: color_data = 12'he21;
			{8'd98, 8'd15}: color_data = 12'he21;
			{8'd98, 8'd16}: color_data = 12'he21;
			{8'd98, 8'd17}: color_data = 12'hf21;
			{8'd98, 8'd18}: color_data = 12'he21;
			{8'd98, 8'd19}: color_data = 12'h500;
			{8'd98, 8'd20}: color_data = 12'h000;
			{8'd98, 8'd21}: color_data = 12'h000;
			{8'd98, 8'd22}: color_data = 12'h020;
			{8'd98, 8'd23}: color_data = 12'h010;
			{8'd98, 8'd24}: color_data = 12'h000;
			{8'd98, 8'd25}: color_data = 12'h000;
			{8'd98, 8'd26}: color_data = 12'h000;
			{8'd98, 8'd27}: color_data = 12'h000;
			{8'd98, 8'd28}: color_data = 12'h000;
			{8'd98, 8'd29}: color_data = 12'h000;
			{8'd98, 8'd30}: color_data = 12'h000;
			{8'd98, 8'd31}: color_data = 12'h000;
			{8'd98, 8'd32}: color_data = 12'h000;
			{8'd98, 8'd33}: color_data = 12'h440;
			{8'd98, 8'd34}: color_data = 12'hfd0;
			{8'd98, 8'd35}: color_data = 12'hfd0;
			{8'd98, 8'd36}: color_data = 12'hfc0;
			{8'd98, 8'd37}: color_data = 12'hfc0;
			{8'd98, 8'd38}: color_data = 12'hfc0;
			{8'd98, 8'd39}: color_data = 12'hfc0;
			{8'd98, 8'd40}: color_data = 12'hfc0;
			{8'd98, 8'd41}: color_data = 12'hfc0;
			{8'd98, 8'd42}: color_data = 12'hfd0;
			{8'd98, 8'd43}: color_data = 12'ha80;
			{8'd98, 8'd44}: color_data = 12'h750;
			{8'd98, 8'd45}: color_data = 12'h970;
			{8'd98, 8'd46}: color_data = 12'hb90;
			{8'd98, 8'd47}: color_data = 12'hca0;
			{8'd98, 8'd48}: color_data = 12'heb0;
			{8'd98, 8'd49}: color_data = 12'hfc0;
			{8'd98, 8'd50}: color_data = 12'hfd0;
			{8'd98, 8'd51}: color_data = 12'hfc0;
			{8'd98, 8'd52}: color_data = 12'hfc0;
			{8'd98, 8'd53}: color_data = 12'hfc0;
			{8'd98, 8'd54}: color_data = 12'hfc0;
			{8'd98, 8'd55}: color_data = 12'hfc0;
			{8'd98, 8'd56}: color_data = 12'hfc0;
			{8'd98, 8'd57}: color_data = 12'hfc0;
			{8'd98, 8'd58}: color_data = 12'hfc0;
			{8'd98, 8'd59}: color_data = 12'hfc0;
			{8'd98, 8'd60}: color_data = 12'hfc0;
			{8'd98, 8'd61}: color_data = 12'hfc0;
			{8'd98, 8'd62}: color_data = 12'hfc0;
			{8'd98, 8'd63}: color_data = 12'hfd0;
			{8'd98, 8'd64}: color_data = 12'hfd0;
			{8'd98, 8'd65}: color_data = 12'hb90;
			{8'd98, 8'd66}: color_data = 12'h220;
			{8'd98, 8'd67}: color_data = 12'h000;
			{8'd98, 8'd68}: color_data = 12'h000;
			{8'd98, 8'd69}: color_data = 12'h000;
			{8'd98, 8'd70}: color_data = 12'h000;
			{8'd98, 8'd71}: color_data = 12'h000;
			{8'd98, 8'd72}: color_data = 12'h000;
			{8'd98, 8'd73}: color_data = 12'h000;
			{8'd98, 8'd74}: color_data = 12'h000;
			{8'd98, 8'd75}: color_data = 12'h000;
			{8'd98, 8'd100}: color_data = 12'he00;
			{8'd98, 8'd101}: color_data = 12'hf01;
			{8'd98, 8'd102}: color_data = 12'he00;
			{8'd98, 8'd103}: color_data = 12'he00;
			{8'd98, 8'd104}: color_data = 12'he00;
			{8'd98, 8'd105}: color_data = 12'he00;
			{8'd98, 8'd106}: color_data = 12'hc00;
			{8'd98, 8'd118}: color_data = 12'he00;
			{8'd98, 8'd119}: color_data = 12'he00;
			{8'd98, 8'd120}: color_data = 12'he00;
			{8'd98, 8'd121}: color_data = 12'he00;
			{8'd98, 8'd122}: color_data = 12'he00;
			{8'd98, 8'd123}: color_data = 12'he00;
			{8'd98, 8'd124}: color_data = 12'he00;
			{8'd98, 8'd125}: color_data = 12'he00;
			{8'd98, 8'd126}: color_data = 12'he00;
			{8'd98, 8'd127}: color_data = 12'he00;
			{8'd98, 8'd128}: color_data = 12'he00;
			{8'd98, 8'd129}: color_data = 12'he00;
			{8'd98, 8'd130}: color_data = 12'he00;
			{8'd98, 8'd131}: color_data = 12'he00;
			{8'd98, 8'd132}: color_data = 12'hf01;
			{8'd98, 8'd133}: color_data = 12'he00;
			{8'd98, 8'd138}: color_data = 12'he00;
			{8'd98, 8'd139}: color_data = 12'he00;
			{8'd98, 8'd140}: color_data = 12'he00;
			{8'd98, 8'd141}: color_data = 12'he00;
			{8'd98, 8'd142}: color_data = 12'he00;
			{8'd98, 8'd143}: color_data = 12'he01;
			{8'd98, 8'd144}: color_data = 12'he00;
			{8'd99, 8'd5}: color_data = 12'h000;
			{8'd99, 8'd6}: color_data = 12'h000;
			{8'd99, 8'd7}: color_data = 12'h000;
			{8'd99, 8'd8}: color_data = 12'h710;
			{8'd99, 8'd9}: color_data = 12'hf21;
			{8'd99, 8'd10}: color_data = 12'he21;
			{8'd99, 8'd11}: color_data = 12'he21;
			{8'd99, 8'd12}: color_data = 12'he21;
			{8'd99, 8'd13}: color_data = 12'he21;
			{8'd99, 8'd14}: color_data = 12'hd20;
			{8'd99, 8'd15}: color_data = 12'hc10;
			{8'd99, 8'd16}: color_data = 12'ha10;
			{8'd99, 8'd17}: color_data = 12'h810;
			{8'd99, 8'd18}: color_data = 12'h400;
			{8'd99, 8'd19}: color_data = 12'h000;
			{8'd99, 8'd20}: color_data = 12'h000;
			{8'd99, 8'd21}: color_data = 12'h251;
			{8'd99, 8'd22}: color_data = 12'h4a3;
			{8'd99, 8'd23}: color_data = 12'h4a3;
			{8'd99, 8'd24}: color_data = 12'h392;
			{8'd99, 8'd25}: color_data = 12'h272;
			{8'd99, 8'd26}: color_data = 12'h251;
			{8'd99, 8'd27}: color_data = 12'h141;
			{8'd99, 8'd28}: color_data = 12'h120;
			{8'd99, 8'd29}: color_data = 12'h010;
			{8'd99, 8'd30}: color_data = 12'h000;
			{8'd99, 8'd31}: color_data = 12'h000;
			{8'd99, 8'd32}: color_data = 12'h000;
			{8'd99, 8'd33}: color_data = 12'h000;
			{8'd99, 8'd34}: color_data = 12'ha80;
			{8'd99, 8'd35}: color_data = 12'hfd0;
			{8'd99, 8'd36}: color_data = 12'hfc0;
			{8'd99, 8'd37}: color_data = 12'hfc0;
			{8'd99, 8'd38}: color_data = 12'hfc0;
			{8'd99, 8'd39}: color_data = 12'hfc0;
			{8'd99, 8'd40}: color_data = 12'hfc0;
			{8'd99, 8'd41}: color_data = 12'hfc0;
			{8'd99, 8'd42}: color_data = 12'hfc0;
			{8'd99, 8'd43}: color_data = 12'hfd0;
			{8'd99, 8'd44}: color_data = 12'hfd0;
			{8'd99, 8'd45}: color_data = 12'hfd0;
			{8'd99, 8'd46}: color_data = 12'hfd0;
			{8'd99, 8'd47}: color_data = 12'hfd0;
			{8'd99, 8'd48}: color_data = 12'hfd0;
			{8'd99, 8'd49}: color_data = 12'hfd0;
			{8'd99, 8'd50}: color_data = 12'hfc0;
			{8'd99, 8'd51}: color_data = 12'hfc0;
			{8'd99, 8'd52}: color_data = 12'hfc0;
			{8'd99, 8'd53}: color_data = 12'hfc0;
			{8'd99, 8'd54}: color_data = 12'hfc0;
			{8'd99, 8'd55}: color_data = 12'hfc0;
			{8'd99, 8'd56}: color_data = 12'hfc0;
			{8'd99, 8'd57}: color_data = 12'hfc0;
			{8'd99, 8'd58}: color_data = 12'hfc0;
			{8'd99, 8'd59}: color_data = 12'hfc0;
			{8'd99, 8'd60}: color_data = 12'hfc0;
			{8'd99, 8'd61}: color_data = 12'hfc0;
			{8'd99, 8'd62}: color_data = 12'hfc0;
			{8'd99, 8'd63}: color_data = 12'hfc0;
			{8'd99, 8'd64}: color_data = 12'hfc0;
			{8'd99, 8'd65}: color_data = 12'hfd0;
			{8'd99, 8'd66}: color_data = 12'hec0;
			{8'd99, 8'd67}: color_data = 12'h750;
			{8'd99, 8'd68}: color_data = 12'h000;
			{8'd99, 8'd69}: color_data = 12'h000;
			{8'd99, 8'd70}: color_data = 12'h000;
			{8'd99, 8'd71}: color_data = 12'h000;
			{8'd99, 8'd72}: color_data = 12'h000;
			{8'd99, 8'd73}: color_data = 12'h000;
			{8'd99, 8'd74}: color_data = 12'h000;
			{8'd99, 8'd75}: color_data = 12'h000;
			{8'd99, 8'd100}: color_data = 12'he00;
			{8'd99, 8'd101}: color_data = 12'hf01;
			{8'd99, 8'd102}: color_data = 12'he00;
			{8'd99, 8'd103}: color_data = 12'he00;
			{8'd99, 8'd104}: color_data = 12'he00;
			{8'd99, 8'd105}: color_data = 12'he00;
			{8'd99, 8'd106}: color_data = 12'hc00;
			{8'd99, 8'd119}: color_data = 12'he00;
			{8'd99, 8'd120}: color_data = 12'he00;
			{8'd99, 8'd121}: color_data = 12'he00;
			{8'd99, 8'd122}: color_data = 12'he01;
			{8'd99, 8'd123}: color_data = 12'he01;
			{8'd99, 8'd124}: color_data = 12'he01;
			{8'd99, 8'd125}: color_data = 12'he01;
			{8'd99, 8'd126}: color_data = 12'he01;
			{8'd99, 8'd127}: color_data = 12'he01;
			{8'd99, 8'd128}: color_data = 12'he01;
			{8'd99, 8'd129}: color_data = 12'he01;
			{8'd99, 8'd130}: color_data = 12'he01;
			{8'd99, 8'd131}: color_data = 12'he01;
			{8'd99, 8'd132}: color_data = 12'hf01;
			{8'd99, 8'd133}: color_data = 12'he00;
			{8'd99, 8'd138}: color_data = 12'he00;
			{8'd99, 8'd139}: color_data = 12'he00;
			{8'd99, 8'd140}: color_data = 12'he00;
			{8'd99, 8'd141}: color_data = 12'he00;
			{8'd99, 8'd142}: color_data = 12'he00;
			{8'd99, 8'd143}: color_data = 12'he01;
			{8'd99, 8'd144}: color_data = 12'he00;
			{8'd100, 8'd2}: color_data = 12'h000;
			{8'd100, 8'd3}: color_data = 12'h000;
			{8'd100, 8'd4}: color_data = 12'h000;
			{8'd100, 8'd5}: color_data = 12'h000;
			{8'd100, 8'd6}: color_data = 12'h000;
			{8'd100, 8'd7}: color_data = 12'h000;
			{8'd100, 8'd8}: color_data = 12'h100;
			{8'd100, 8'd9}: color_data = 12'h910;
			{8'd100, 8'd10}: color_data = 12'h910;
			{8'd100, 8'd11}: color_data = 12'h710;
			{8'd100, 8'd12}: color_data = 12'h500;
			{8'd100, 8'd13}: color_data = 12'h300;
			{8'd100, 8'd14}: color_data = 12'h100;
			{8'd100, 8'd15}: color_data = 12'h000;
			{8'd100, 8'd16}: color_data = 12'h000;
			{8'd100, 8'd17}: color_data = 12'h000;
			{8'd100, 8'd18}: color_data = 12'h000;
			{8'd100, 8'd19}: color_data = 12'h000;
			{8'd100, 8'd20}: color_data = 12'h141;
			{8'd100, 8'd21}: color_data = 12'h4b3;
			{8'd100, 8'd22}: color_data = 12'h4b3;
			{8'd100, 8'd23}: color_data = 12'h4b3;
			{8'd100, 8'd24}: color_data = 12'h4b3;
			{8'd100, 8'd25}: color_data = 12'h4b3;
			{8'd100, 8'd26}: color_data = 12'h4b3;
			{8'd100, 8'd27}: color_data = 12'h4b3;
			{8'd100, 8'd28}: color_data = 12'h4b3;
			{8'd100, 8'd29}: color_data = 12'h372;
			{8'd100, 8'd30}: color_data = 12'h000;
			{8'd100, 8'd31}: color_data = 12'h000;
			{8'd100, 8'd32}: color_data = 12'h000;
			{8'd100, 8'd33}: color_data = 12'h000;
			{8'd100, 8'd34}: color_data = 12'h220;
			{8'd100, 8'd35}: color_data = 12'hfc0;
			{8'd100, 8'd36}: color_data = 12'hfd0;
			{8'd100, 8'd37}: color_data = 12'hfc0;
			{8'd100, 8'd38}: color_data = 12'hfc0;
			{8'd100, 8'd39}: color_data = 12'hfc0;
			{8'd100, 8'd40}: color_data = 12'hfc0;
			{8'd100, 8'd41}: color_data = 12'hfc0;
			{8'd100, 8'd42}: color_data = 12'hfc0;
			{8'd100, 8'd43}: color_data = 12'hfc0;
			{8'd100, 8'd44}: color_data = 12'hfc0;
			{8'd100, 8'd45}: color_data = 12'hfc0;
			{8'd100, 8'd46}: color_data = 12'hfc0;
			{8'd100, 8'd47}: color_data = 12'hfc0;
			{8'd100, 8'd48}: color_data = 12'hfc0;
			{8'd100, 8'd49}: color_data = 12'hfc0;
			{8'd100, 8'd50}: color_data = 12'hfc0;
			{8'd100, 8'd51}: color_data = 12'hfc0;
			{8'd100, 8'd52}: color_data = 12'hfc0;
			{8'd100, 8'd53}: color_data = 12'hfc0;
			{8'd100, 8'd54}: color_data = 12'hfc0;
			{8'd100, 8'd55}: color_data = 12'hfd0;
			{8'd100, 8'd56}: color_data = 12'hfd0;
			{8'd100, 8'd57}: color_data = 12'hfc0;
			{8'd100, 8'd58}: color_data = 12'hfc0;
			{8'd100, 8'd59}: color_data = 12'hfc0;
			{8'd100, 8'd60}: color_data = 12'hfc0;
			{8'd100, 8'd61}: color_data = 12'hfc0;
			{8'd100, 8'd62}: color_data = 12'hfc0;
			{8'd100, 8'd63}: color_data = 12'hfc0;
			{8'd100, 8'd64}: color_data = 12'hfc0;
			{8'd100, 8'd65}: color_data = 12'hfc0;
			{8'd100, 8'd66}: color_data = 12'hfd0;
			{8'd100, 8'd67}: color_data = 12'hec0;
			{8'd100, 8'd68}: color_data = 12'h210;
			{8'd100, 8'd69}: color_data = 12'h000;
			{8'd100, 8'd70}: color_data = 12'h000;
			{8'd100, 8'd71}: color_data = 12'h000;
			{8'd100, 8'd72}: color_data = 12'h000;
			{8'd100, 8'd73}: color_data = 12'h000;
			{8'd100, 8'd74}: color_data = 12'h000;
			{8'd100, 8'd75}: color_data = 12'h000;
			{8'd100, 8'd100}: color_data = 12'he00;
			{8'd100, 8'd101}: color_data = 12'hf01;
			{8'd100, 8'd102}: color_data = 12'he00;
			{8'd100, 8'd103}: color_data = 12'he00;
			{8'd100, 8'd104}: color_data = 12'he00;
			{8'd100, 8'd105}: color_data = 12'he00;
			{8'd100, 8'd106}: color_data = 12'hc00;
			{8'd100, 8'd120}: color_data = 12'hd00;
			{8'd100, 8'd121}: color_data = 12'he01;
			{8'd100, 8'd122}: color_data = 12'he00;
			{8'd100, 8'd123}: color_data = 12'he00;
			{8'd100, 8'd124}: color_data = 12'he00;
			{8'd100, 8'd125}: color_data = 12'he00;
			{8'd100, 8'd126}: color_data = 12'he00;
			{8'd100, 8'd127}: color_data = 12'he00;
			{8'd100, 8'd128}: color_data = 12'he00;
			{8'd100, 8'd129}: color_data = 12'he00;
			{8'd100, 8'd130}: color_data = 12'he00;
			{8'd100, 8'd131}: color_data = 12'he00;
			{8'd100, 8'd132}: color_data = 12'he00;
			{8'd100, 8'd133}: color_data = 12'he00;
			{8'd100, 8'd138}: color_data = 12'he00;
			{8'd100, 8'd139}: color_data = 12'he00;
			{8'd100, 8'd140}: color_data = 12'he00;
			{8'd100, 8'd141}: color_data = 12'he00;
			{8'd100, 8'd142}: color_data = 12'he00;
			{8'd100, 8'd143}: color_data = 12'he01;
			{8'd100, 8'd144}: color_data = 12'he00;
			{8'd101, 8'd2}: color_data = 12'h000;
			{8'd101, 8'd3}: color_data = 12'h000;
			{8'd101, 8'd4}: color_data = 12'h000;
			{8'd101, 8'd5}: color_data = 12'h000;
			{8'd101, 8'd6}: color_data = 12'h000;
			{8'd101, 8'd7}: color_data = 12'h000;
			{8'd101, 8'd8}: color_data = 12'h000;
			{8'd101, 8'd9}: color_data = 12'h000;
			{8'd101, 8'd10}: color_data = 12'h000;
			{8'd101, 8'd11}: color_data = 12'h000;
			{8'd101, 8'd12}: color_data = 12'h000;
			{8'd101, 8'd13}: color_data = 12'h000;
			{8'd101, 8'd14}: color_data = 12'h000;
			{8'd101, 8'd15}: color_data = 12'h000;
			{8'd101, 8'd16}: color_data = 12'h000;
			{8'd101, 8'd17}: color_data = 12'h010;
			{8'd101, 8'd18}: color_data = 12'h120;
			{8'd101, 8'd19}: color_data = 12'h251;
			{8'd101, 8'd20}: color_data = 12'h4a3;
			{8'd101, 8'd21}: color_data = 12'h4b3;
			{8'd101, 8'd22}: color_data = 12'h4a3;
			{8'd101, 8'd23}: color_data = 12'h4a3;
			{8'd101, 8'd24}: color_data = 12'h4a3;
			{8'd101, 8'd25}: color_data = 12'h4a3;
			{8'd101, 8'd26}: color_data = 12'h4a3;
			{8'd101, 8'd27}: color_data = 12'h4a3;
			{8'd101, 8'd28}: color_data = 12'h4b3;
			{8'd101, 8'd29}: color_data = 12'h382;
			{8'd101, 8'd30}: color_data = 12'h000;
			{8'd101, 8'd31}: color_data = 12'h000;
			{8'd101, 8'd32}: color_data = 12'h000;
			{8'd101, 8'd33}: color_data = 12'h000;
			{8'd101, 8'd34}: color_data = 12'h000;
			{8'd101, 8'd35}: color_data = 12'h870;
			{8'd101, 8'd36}: color_data = 12'hfd0;
			{8'd101, 8'd37}: color_data = 12'hfc0;
			{8'd101, 8'd38}: color_data = 12'hfc0;
			{8'd101, 8'd39}: color_data = 12'hfc0;
			{8'd101, 8'd40}: color_data = 12'hfc0;
			{8'd101, 8'd41}: color_data = 12'hfc0;
			{8'd101, 8'd42}: color_data = 12'hfc0;
			{8'd101, 8'd43}: color_data = 12'hfc0;
			{8'd101, 8'd44}: color_data = 12'hfc0;
			{8'd101, 8'd45}: color_data = 12'hfc0;
			{8'd101, 8'd46}: color_data = 12'hfc0;
			{8'd101, 8'd47}: color_data = 12'hfc0;
			{8'd101, 8'd48}: color_data = 12'hfc0;
			{8'd101, 8'd49}: color_data = 12'hfc0;
			{8'd101, 8'd50}: color_data = 12'hfc0;
			{8'd101, 8'd51}: color_data = 12'hfc0;
			{8'd101, 8'd52}: color_data = 12'hfc0;
			{8'd101, 8'd53}: color_data = 12'hfc0;
			{8'd101, 8'd54}: color_data = 12'hfd0;
			{8'd101, 8'd55}: color_data = 12'hb90;
			{8'd101, 8'd56}: color_data = 12'hfc0;
			{8'd101, 8'd57}: color_data = 12'hfd0;
			{8'd101, 8'd58}: color_data = 12'hfc0;
			{8'd101, 8'd59}: color_data = 12'hfc0;
			{8'd101, 8'd60}: color_data = 12'hfc0;
			{8'd101, 8'd61}: color_data = 12'hfc0;
			{8'd101, 8'd62}: color_data = 12'hfc0;
			{8'd101, 8'd63}: color_data = 12'hfc0;
			{8'd101, 8'd64}: color_data = 12'hfc0;
			{8'd101, 8'd65}: color_data = 12'hfc0;
			{8'd101, 8'd66}: color_data = 12'hfd0;
			{8'd101, 8'd67}: color_data = 12'ha80;
			{8'd101, 8'd68}: color_data = 12'h000;
			{8'd101, 8'd69}: color_data = 12'h000;
			{8'd101, 8'd70}: color_data = 12'h000;
			{8'd101, 8'd71}: color_data = 12'h000;
			{8'd101, 8'd72}: color_data = 12'h000;
			{8'd101, 8'd73}: color_data = 12'h000;
			{8'd101, 8'd74}: color_data = 12'h000;
			{8'd101, 8'd100}: color_data = 12'he00;
			{8'd101, 8'd101}: color_data = 12'hf01;
			{8'd101, 8'd102}: color_data = 12'he00;
			{8'd101, 8'd103}: color_data = 12'he00;
			{8'd101, 8'd104}: color_data = 12'he00;
			{8'd101, 8'd105}: color_data = 12'he00;
			{8'd101, 8'd106}: color_data = 12'hc00;
			{8'd101, 8'd132}: color_data = 12'hf00;
			{8'd101, 8'd133}: color_data = 12'he00;
			{8'd101, 8'd138}: color_data = 12'he00;
			{8'd101, 8'd139}: color_data = 12'he00;
			{8'd101, 8'd140}: color_data = 12'he00;
			{8'd101, 8'd141}: color_data = 12'he00;
			{8'd101, 8'd142}: color_data = 12'he00;
			{8'd101, 8'd143}: color_data = 12'he01;
			{8'd101, 8'd144}: color_data = 12'he00;
			{8'd102, 8'd2}: color_data = 12'h000;
			{8'd102, 8'd3}: color_data = 12'h000;
			{8'd102, 8'd4}: color_data = 12'h000;
			{8'd102, 8'd5}: color_data = 12'h262;
			{8'd102, 8'd6}: color_data = 12'h393;
			{8'd102, 8'd7}: color_data = 12'h261;
			{8'd102, 8'd8}: color_data = 12'h000;
			{8'd102, 8'd9}: color_data = 12'h000;
			{8'd102, 8'd10}: color_data = 12'h010;
			{8'd102, 8'd11}: color_data = 12'h120;
			{8'd102, 8'd12}: color_data = 12'h141;
			{8'd102, 8'd13}: color_data = 12'h251;
			{8'd102, 8'd14}: color_data = 12'h272;
			{8'd102, 8'd15}: color_data = 12'h382;
			{8'd102, 8'd16}: color_data = 12'h392;
			{8'd102, 8'd17}: color_data = 12'h4a3;
			{8'd102, 8'd18}: color_data = 12'h4b3;
			{8'd102, 8'd19}: color_data = 12'h4b3;
			{8'd102, 8'd20}: color_data = 12'h4b3;
			{8'd102, 8'd21}: color_data = 12'h4a3;
			{8'd102, 8'd22}: color_data = 12'h4a3;
			{8'd102, 8'd23}: color_data = 12'h4a3;
			{8'd102, 8'd24}: color_data = 12'h4a3;
			{8'd102, 8'd25}: color_data = 12'h4a3;
			{8'd102, 8'd26}: color_data = 12'h4a3;
			{8'd102, 8'd27}: color_data = 12'h4a3;
			{8'd102, 8'd28}: color_data = 12'h4b3;
			{8'd102, 8'd29}: color_data = 12'h382;
			{8'd102, 8'd30}: color_data = 12'h000;
			{8'd102, 8'd31}: color_data = 12'h000;
			{8'd102, 8'd32}: color_data = 12'h000;
			{8'd102, 8'd33}: color_data = 12'h000;
			{8'd102, 8'd34}: color_data = 12'h000;
			{8'd102, 8'd35}: color_data = 12'h110;
			{8'd102, 8'd36}: color_data = 12'hdb0;
			{8'd102, 8'd37}: color_data = 12'hfd0;
			{8'd102, 8'd38}: color_data = 12'hfc0;
			{8'd102, 8'd39}: color_data = 12'hfc0;
			{8'd102, 8'd40}: color_data = 12'hfc0;
			{8'd102, 8'd41}: color_data = 12'hfc0;
			{8'd102, 8'd42}: color_data = 12'hfc0;
			{8'd102, 8'd43}: color_data = 12'hfc0;
			{8'd102, 8'd44}: color_data = 12'hfc0;
			{8'd102, 8'd45}: color_data = 12'hfc0;
			{8'd102, 8'd46}: color_data = 12'hfc0;
			{8'd102, 8'd47}: color_data = 12'hfc0;
			{8'd102, 8'd48}: color_data = 12'hfc0;
			{8'd102, 8'd49}: color_data = 12'hfc0;
			{8'd102, 8'd50}: color_data = 12'hfc0;
			{8'd102, 8'd51}: color_data = 12'hfc0;
			{8'd102, 8'd52}: color_data = 12'hfc0;
			{8'd102, 8'd53}: color_data = 12'hfd0;
			{8'd102, 8'd54}: color_data = 12'hca0;
			{8'd102, 8'd55}: color_data = 12'h000;
			{8'd102, 8'd56}: color_data = 12'h870;
			{8'd102, 8'd57}: color_data = 12'hfd0;
			{8'd102, 8'd58}: color_data = 12'hfc0;
			{8'd102, 8'd59}: color_data = 12'hfc0;
			{8'd102, 8'd60}: color_data = 12'hfc0;
			{8'd102, 8'd61}: color_data = 12'hfc0;
			{8'd102, 8'd62}: color_data = 12'hfc0;
			{8'd102, 8'd63}: color_data = 12'hfc0;
			{8'd102, 8'd64}: color_data = 12'hfc0;
			{8'd102, 8'd65}: color_data = 12'hfd0;
			{8'd102, 8'd66}: color_data = 12'hfd0;
			{8'd102, 8'd67}: color_data = 12'h430;
			{8'd102, 8'd68}: color_data = 12'h000;
			{8'd102, 8'd69}: color_data = 12'h000;
			{8'd102, 8'd70}: color_data = 12'h000;
			{8'd102, 8'd71}: color_data = 12'h000;
			{8'd102, 8'd72}: color_data = 12'h000;
			{8'd102, 8'd73}: color_data = 12'h000;
			{8'd102, 8'd74}: color_data = 12'h000;
			{8'd102, 8'd100}: color_data = 12'he00;
			{8'd102, 8'd101}: color_data = 12'hf01;
			{8'd102, 8'd102}: color_data = 12'he00;
			{8'd102, 8'd103}: color_data = 12'he00;
			{8'd102, 8'd104}: color_data = 12'he00;
			{8'd102, 8'd105}: color_data = 12'he00;
			{8'd102, 8'd106}: color_data = 12'hc00;
			{8'd102, 8'd138}: color_data = 12'he00;
			{8'd102, 8'd139}: color_data = 12'he00;
			{8'd102, 8'd140}: color_data = 12'he00;
			{8'd102, 8'd141}: color_data = 12'he00;
			{8'd102, 8'd142}: color_data = 12'he00;
			{8'd102, 8'd143}: color_data = 12'he01;
			{8'd102, 8'd144}: color_data = 12'he00;
			{8'd103, 8'd2}: color_data = 12'h000;
			{8'd103, 8'd3}: color_data = 12'h000;
			{8'd103, 8'd4}: color_data = 12'h010;
			{8'd103, 8'd5}: color_data = 12'h4a3;
			{8'd103, 8'd6}: color_data = 12'h4b3;
			{8'd103, 8'd7}: color_data = 12'h4a3;
			{8'd103, 8'd8}: color_data = 12'h382;
			{8'd103, 8'd9}: color_data = 12'h392;
			{8'd103, 8'd10}: color_data = 12'h4a3;
			{8'd103, 8'd11}: color_data = 12'h4b3;
			{8'd103, 8'd12}: color_data = 12'h4b3;
			{8'd103, 8'd13}: color_data = 12'h4b3;
			{8'd103, 8'd14}: color_data = 12'h4b3;
			{8'd103, 8'd15}: color_data = 12'h4b3;
			{8'd103, 8'd16}: color_data = 12'h4b3;
			{8'd103, 8'd17}: color_data = 12'h4b3;
			{8'd103, 8'd18}: color_data = 12'h4a3;
			{8'd103, 8'd19}: color_data = 12'h4a3;
			{8'd103, 8'd20}: color_data = 12'h4a3;
			{8'd103, 8'd21}: color_data = 12'h4a3;
			{8'd103, 8'd22}: color_data = 12'h4a3;
			{8'd103, 8'd23}: color_data = 12'h4a3;
			{8'd103, 8'd24}: color_data = 12'h4a3;
			{8'd103, 8'd25}: color_data = 12'h4a3;
			{8'd103, 8'd26}: color_data = 12'h4a3;
			{8'd103, 8'd27}: color_data = 12'h4a3;
			{8'd103, 8'd28}: color_data = 12'h4b3;
			{8'd103, 8'd29}: color_data = 12'h392;
			{8'd103, 8'd30}: color_data = 12'h000;
			{8'd103, 8'd31}: color_data = 12'h000;
			{8'd103, 8'd32}: color_data = 12'h000;
			{8'd103, 8'd33}: color_data = 12'h000;
			{8'd103, 8'd34}: color_data = 12'h000;
			{8'd103, 8'd35}: color_data = 12'h000;
			{8'd103, 8'd36}: color_data = 12'h650;
			{8'd103, 8'd37}: color_data = 12'hfd0;
			{8'd103, 8'd38}: color_data = 12'hfc0;
			{8'd103, 8'd39}: color_data = 12'hfc0;
			{8'd103, 8'd40}: color_data = 12'hfc0;
			{8'd103, 8'd41}: color_data = 12'hfc0;
			{8'd103, 8'd42}: color_data = 12'hfc0;
			{8'd103, 8'd43}: color_data = 12'hfc0;
			{8'd103, 8'd44}: color_data = 12'hfc0;
			{8'd103, 8'd45}: color_data = 12'hfc0;
			{8'd103, 8'd46}: color_data = 12'hfc0;
			{8'd103, 8'd47}: color_data = 12'hfc0;
			{8'd103, 8'd48}: color_data = 12'hfc0;
			{8'd103, 8'd49}: color_data = 12'hfc0;
			{8'd103, 8'd50}: color_data = 12'hfc0;
			{8'd103, 8'd51}: color_data = 12'hfc0;
			{8'd103, 8'd52}: color_data = 12'hfd0;
			{8'd103, 8'd53}: color_data = 12'hfd0;
			{8'd103, 8'd54}: color_data = 12'h540;
			{8'd103, 8'd55}: color_data = 12'h000;
			{8'd103, 8'd56}: color_data = 12'h000;
			{8'd103, 8'd57}: color_data = 12'hb90;
			{8'd103, 8'd58}: color_data = 12'hfd0;
			{8'd103, 8'd59}: color_data = 12'hfc0;
			{8'd103, 8'd60}: color_data = 12'hfc0;
			{8'd103, 8'd61}: color_data = 12'hfc0;
			{8'd103, 8'd62}: color_data = 12'hfc0;
			{8'd103, 8'd63}: color_data = 12'hfc0;
			{8'd103, 8'd64}: color_data = 12'hfc0;
			{8'd103, 8'd65}: color_data = 12'hfd0;
			{8'd103, 8'd66}: color_data = 12'hb90;
			{8'd103, 8'd67}: color_data = 12'h000;
			{8'd103, 8'd68}: color_data = 12'h000;
			{8'd103, 8'd69}: color_data = 12'h000;
			{8'd103, 8'd70}: color_data = 12'h000;
			{8'd103, 8'd71}: color_data = 12'h000;
			{8'd103, 8'd72}: color_data = 12'h000;
			{8'd103, 8'd73}: color_data = 12'h000;
			{8'd103, 8'd74}: color_data = 12'h000;
			{8'd103, 8'd100}: color_data = 12'he00;
			{8'd103, 8'd101}: color_data = 12'hf01;
			{8'd103, 8'd102}: color_data = 12'he00;
			{8'd103, 8'd103}: color_data = 12'he00;
			{8'd103, 8'd104}: color_data = 12'he00;
			{8'd103, 8'd105}: color_data = 12'he00;
			{8'd103, 8'd106}: color_data = 12'hc00;
			{8'd103, 8'd121}: color_data = 12'hd00;
			{8'd103, 8'd122}: color_data = 12'he00;
			{8'd103, 8'd123}: color_data = 12'he00;
			{8'd103, 8'd124}: color_data = 12'he00;
			{8'd103, 8'd125}: color_data = 12'he00;
			{8'd103, 8'd126}: color_data = 12'he00;
			{8'd103, 8'd127}: color_data = 12'he00;
			{8'd103, 8'd128}: color_data = 12'he00;
			{8'd103, 8'd129}: color_data = 12'hd00;
			{8'd103, 8'd138}: color_data = 12'he00;
			{8'd103, 8'd139}: color_data = 12'he00;
			{8'd103, 8'd140}: color_data = 12'he00;
			{8'd103, 8'd141}: color_data = 12'he00;
			{8'd103, 8'd142}: color_data = 12'he00;
			{8'd103, 8'd143}: color_data = 12'he01;
			{8'd103, 8'd144}: color_data = 12'he00;
			{8'd104, 8'd2}: color_data = 12'h000;
			{8'd104, 8'd3}: color_data = 12'h000;
			{8'd104, 8'd4}: color_data = 12'h000;
			{8'd104, 8'd5}: color_data = 12'h382;
			{8'd104, 8'd6}: color_data = 12'h4b3;
			{8'd104, 8'd7}: color_data = 12'h4b3;
			{8'd104, 8'd8}: color_data = 12'h4b3;
			{8'd104, 8'd9}: color_data = 12'h4b3;
			{8'd104, 8'd10}: color_data = 12'h4b3;
			{8'd104, 8'd11}: color_data = 12'h4b3;
			{8'd104, 8'd12}: color_data = 12'h4a3;
			{8'd104, 8'd13}: color_data = 12'h4a3;
			{8'd104, 8'd14}: color_data = 12'h4a3;
			{8'd104, 8'd15}: color_data = 12'h4a3;
			{8'd104, 8'd16}: color_data = 12'h4a3;
			{8'd104, 8'd17}: color_data = 12'h4a3;
			{8'd104, 8'd18}: color_data = 12'h4a3;
			{8'd104, 8'd19}: color_data = 12'h4a3;
			{8'd104, 8'd20}: color_data = 12'h4a3;
			{8'd104, 8'd21}: color_data = 12'h4a3;
			{8'd104, 8'd22}: color_data = 12'h4a3;
			{8'd104, 8'd23}: color_data = 12'h4a3;
			{8'd104, 8'd24}: color_data = 12'h4a3;
			{8'd104, 8'd25}: color_data = 12'h4a3;
			{8'd104, 8'd26}: color_data = 12'h4a3;
			{8'd104, 8'd27}: color_data = 12'h4a3;
			{8'd104, 8'd28}: color_data = 12'h4b3;
			{8'd104, 8'd29}: color_data = 12'h392;
			{8'd104, 8'd30}: color_data = 12'h000;
			{8'd104, 8'd31}: color_data = 12'h000;
			{8'd104, 8'd32}: color_data = 12'h000;
			{8'd104, 8'd33}: color_data = 12'h000;
			{8'd104, 8'd34}: color_data = 12'h000;
			{8'd104, 8'd35}: color_data = 12'h000;
			{8'd104, 8'd36}: color_data = 12'h000;
			{8'd104, 8'd37}: color_data = 12'hb90;
			{8'd104, 8'd38}: color_data = 12'hfd0;
			{8'd104, 8'd39}: color_data = 12'hfc0;
			{8'd104, 8'd40}: color_data = 12'hfc0;
			{8'd104, 8'd41}: color_data = 12'hfc0;
			{8'd104, 8'd42}: color_data = 12'hfc0;
			{8'd104, 8'd43}: color_data = 12'hfc0;
			{8'd104, 8'd44}: color_data = 12'hfc0;
			{8'd104, 8'd45}: color_data = 12'hfc0;
			{8'd104, 8'd46}: color_data = 12'hfc0;
			{8'd104, 8'd47}: color_data = 12'hfc0;
			{8'd104, 8'd48}: color_data = 12'hfc0;
			{8'd104, 8'd49}: color_data = 12'hfc0;
			{8'd104, 8'd50}: color_data = 12'hfc0;
			{8'd104, 8'd51}: color_data = 12'hfc0;
			{8'd104, 8'd52}: color_data = 12'hfd0;
			{8'd104, 8'd53}: color_data = 12'ha90;
			{8'd104, 8'd54}: color_data = 12'h000;
			{8'd104, 8'd55}: color_data = 12'h000;
			{8'd104, 8'd56}: color_data = 12'h000;
			{8'd104, 8'd57}: color_data = 12'h110;
			{8'd104, 8'd58}: color_data = 12'hda0;
			{8'd104, 8'd59}: color_data = 12'hfd0;
			{8'd104, 8'd60}: color_data = 12'hfc0;
			{8'd104, 8'd61}: color_data = 12'hfc0;
			{8'd104, 8'd62}: color_data = 12'hfc0;
			{8'd104, 8'd63}: color_data = 12'hfc0;
			{8'd104, 8'd64}: color_data = 12'hfc0;
			{8'd104, 8'd65}: color_data = 12'hfd0;
			{8'd104, 8'd66}: color_data = 12'h540;
			{8'd104, 8'd67}: color_data = 12'h000;
			{8'd104, 8'd68}: color_data = 12'h000;
			{8'd104, 8'd69}: color_data = 12'h000;
			{8'd104, 8'd70}: color_data = 12'h000;
			{8'd104, 8'd71}: color_data = 12'h000;
			{8'd104, 8'd72}: color_data = 12'h000;
			{8'd104, 8'd73}: color_data = 12'h000;
			{8'd104, 8'd100}: color_data = 12'he00;
			{8'd104, 8'd101}: color_data = 12'hf01;
			{8'd104, 8'd102}: color_data = 12'he00;
			{8'd104, 8'd103}: color_data = 12'he00;
			{8'd104, 8'd104}: color_data = 12'he00;
			{8'd104, 8'd105}: color_data = 12'he00;
			{8'd104, 8'd106}: color_data = 12'hc00;
			{8'd104, 8'd119}: color_data = 12'hf00;
			{8'd104, 8'd120}: color_data = 12'he00;
			{8'd104, 8'd121}: color_data = 12'he00;
			{8'd104, 8'd122}: color_data = 12'he00;
			{8'd104, 8'd123}: color_data = 12'he01;
			{8'd104, 8'd124}: color_data = 12'hf01;
			{8'd104, 8'd125}: color_data = 12'he01;
			{8'd104, 8'd126}: color_data = 12'hf01;
			{8'd104, 8'd127}: color_data = 12'he01;
			{8'd104, 8'd128}: color_data = 12'he00;
			{8'd104, 8'd129}: color_data = 12'he00;
			{8'd104, 8'd130}: color_data = 12'he00;
			{8'd104, 8'd131}: color_data = 12'hf01;
			{8'd104, 8'd138}: color_data = 12'he00;
			{8'd104, 8'd139}: color_data = 12'he00;
			{8'd104, 8'd140}: color_data = 12'he00;
			{8'd104, 8'd141}: color_data = 12'he00;
			{8'd104, 8'd142}: color_data = 12'he00;
			{8'd104, 8'd143}: color_data = 12'he01;
			{8'd104, 8'd144}: color_data = 12'he00;
			{8'd105, 8'd2}: color_data = 12'h000;
			{8'd105, 8'd3}: color_data = 12'h000;
			{8'd105, 8'd4}: color_data = 12'h000;
			{8'd105, 8'd5}: color_data = 12'h272;
			{8'd105, 8'd6}: color_data = 12'h4b3;
			{8'd105, 8'd7}: color_data = 12'h4a3;
			{8'd105, 8'd8}: color_data = 12'h4a3;
			{8'd105, 8'd9}: color_data = 12'h4a3;
			{8'd105, 8'd10}: color_data = 12'h4a3;
			{8'd105, 8'd11}: color_data = 12'h4a3;
			{8'd105, 8'd12}: color_data = 12'h4a3;
			{8'd105, 8'd13}: color_data = 12'h4a3;
			{8'd105, 8'd14}: color_data = 12'h4a3;
			{8'd105, 8'd15}: color_data = 12'h4a3;
			{8'd105, 8'd16}: color_data = 12'h4a3;
			{8'd105, 8'd17}: color_data = 12'h4a3;
			{8'd105, 8'd18}: color_data = 12'h4a3;
			{8'd105, 8'd19}: color_data = 12'h4a3;
			{8'd105, 8'd20}: color_data = 12'h4a3;
			{8'd105, 8'd21}: color_data = 12'h4a3;
			{8'd105, 8'd22}: color_data = 12'h4a3;
			{8'd105, 8'd23}: color_data = 12'h4a3;
			{8'd105, 8'd24}: color_data = 12'h4a3;
			{8'd105, 8'd25}: color_data = 12'h4a3;
			{8'd105, 8'd26}: color_data = 12'h4a3;
			{8'd105, 8'd27}: color_data = 12'h4a3;
			{8'd105, 8'd28}: color_data = 12'h4b3;
			{8'd105, 8'd29}: color_data = 12'h392;
			{8'd105, 8'd30}: color_data = 12'h000;
			{8'd105, 8'd31}: color_data = 12'h000;
			{8'd105, 8'd32}: color_data = 12'h000;
			{8'd105, 8'd33}: color_data = 12'h000;
			{8'd105, 8'd34}: color_data = 12'h000;
			{8'd105, 8'd35}: color_data = 12'h000;
			{8'd105, 8'd36}: color_data = 12'h000;
			{8'd105, 8'd37}: color_data = 12'h330;
			{8'd105, 8'd38}: color_data = 12'hfc0;
			{8'd105, 8'd39}: color_data = 12'hfd0;
			{8'd105, 8'd40}: color_data = 12'hfc0;
			{8'd105, 8'd41}: color_data = 12'hfc0;
			{8'd105, 8'd42}: color_data = 12'hfc0;
			{8'd105, 8'd43}: color_data = 12'hfc0;
			{8'd105, 8'd44}: color_data = 12'hfc0;
			{8'd105, 8'd45}: color_data = 12'hfc0;
			{8'd105, 8'd46}: color_data = 12'hfc0;
			{8'd105, 8'd47}: color_data = 12'hfc0;
			{8'd105, 8'd48}: color_data = 12'hfc0;
			{8'd105, 8'd49}: color_data = 12'hfc0;
			{8'd105, 8'd50}: color_data = 12'hfc0;
			{8'd105, 8'd51}: color_data = 12'hfd0;
			{8'd105, 8'd52}: color_data = 12'hfc0;
			{8'd105, 8'd53}: color_data = 12'h220;
			{8'd105, 8'd54}: color_data = 12'h000;
			{8'd105, 8'd55}: color_data = 12'h000;
			{8'd105, 8'd56}: color_data = 12'h000;
			{8'd105, 8'd57}: color_data = 12'h000;
			{8'd105, 8'd58}: color_data = 12'h320;
			{8'd105, 8'd59}: color_data = 12'hec0;
			{8'd105, 8'd60}: color_data = 12'hfd0;
			{8'd105, 8'd61}: color_data = 12'hfc0;
			{8'd105, 8'd62}: color_data = 12'hfc0;
			{8'd105, 8'd63}: color_data = 12'hfc0;
			{8'd105, 8'd64}: color_data = 12'hfd0;
			{8'd105, 8'd65}: color_data = 12'hda0;
			{8'd105, 8'd66}: color_data = 12'h000;
			{8'd105, 8'd67}: color_data = 12'h000;
			{8'd105, 8'd68}: color_data = 12'h000;
			{8'd105, 8'd69}: color_data = 12'h000;
			{8'd105, 8'd70}: color_data = 12'h000;
			{8'd105, 8'd71}: color_data = 12'h000;
			{8'd105, 8'd72}: color_data = 12'h000;
			{8'd105, 8'd73}: color_data = 12'h000;
			{8'd105, 8'd100}: color_data = 12'he00;
			{8'd105, 8'd101}: color_data = 12'hf01;
			{8'd105, 8'd102}: color_data = 12'he00;
			{8'd105, 8'd103}: color_data = 12'he00;
			{8'd105, 8'd104}: color_data = 12'he00;
			{8'd105, 8'd105}: color_data = 12'he00;
			{8'd105, 8'd106}: color_data = 12'hc00;
			{8'd105, 8'd118}: color_data = 12'hf00;
			{8'd105, 8'd119}: color_data = 12'he00;
			{8'd105, 8'd120}: color_data = 12'he01;
			{8'd105, 8'd121}: color_data = 12'he00;
			{8'd105, 8'd122}: color_data = 12'he00;
			{8'd105, 8'd123}: color_data = 12'he00;
			{8'd105, 8'd124}: color_data = 12'he00;
			{8'd105, 8'd125}: color_data = 12'he00;
			{8'd105, 8'd126}: color_data = 12'he00;
			{8'd105, 8'd127}: color_data = 12'he00;
			{8'd105, 8'd128}: color_data = 12'he00;
			{8'd105, 8'd129}: color_data = 12'he00;
			{8'd105, 8'd130}: color_data = 12'he01;
			{8'd105, 8'd131}: color_data = 12'he00;
			{8'd105, 8'd132}: color_data = 12'he00;
			{8'd105, 8'd138}: color_data = 12'he00;
			{8'd105, 8'd139}: color_data = 12'he00;
			{8'd105, 8'd140}: color_data = 12'he00;
			{8'd105, 8'd141}: color_data = 12'he00;
			{8'd105, 8'd142}: color_data = 12'he00;
			{8'd105, 8'd143}: color_data = 12'he01;
			{8'd105, 8'd144}: color_data = 12'he00;
			{8'd106, 8'd3}: color_data = 12'h000;
			{8'd106, 8'd4}: color_data = 12'h000;
			{8'd106, 8'd5}: color_data = 12'h251;
			{8'd106, 8'd6}: color_data = 12'h4b3;
			{8'd106, 8'd7}: color_data = 12'h4a3;
			{8'd106, 8'd8}: color_data = 12'h4a3;
			{8'd106, 8'd9}: color_data = 12'h4a3;
			{8'd106, 8'd10}: color_data = 12'h4a3;
			{8'd106, 8'd11}: color_data = 12'h4a3;
			{8'd106, 8'd12}: color_data = 12'h4a3;
			{8'd106, 8'd13}: color_data = 12'h4a3;
			{8'd106, 8'd14}: color_data = 12'h4a3;
			{8'd106, 8'd15}: color_data = 12'h4a3;
			{8'd106, 8'd16}: color_data = 12'h4a3;
			{8'd106, 8'd17}: color_data = 12'h4a3;
			{8'd106, 8'd18}: color_data = 12'h4a3;
			{8'd106, 8'd19}: color_data = 12'h4a3;
			{8'd106, 8'd20}: color_data = 12'h4b3;
			{8'd106, 8'd21}: color_data = 12'h4b3;
			{8'd106, 8'd22}: color_data = 12'h4b3;
			{8'd106, 8'd23}: color_data = 12'h4b3;
			{8'd106, 8'd24}: color_data = 12'h4a3;
			{8'd106, 8'd25}: color_data = 12'h4a3;
			{8'd106, 8'd26}: color_data = 12'h4a3;
			{8'd106, 8'd27}: color_data = 12'h4a3;
			{8'd106, 8'd28}: color_data = 12'h4b3;
			{8'd106, 8'd29}: color_data = 12'h393;
			{8'd106, 8'd30}: color_data = 12'h000;
			{8'd106, 8'd31}: color_data = 12'h000;
			{8'd106, 8'd32}: color_data = 12'h000;
			{8'd106, 8'd33}: color_data = 12'h000;
			{8'd106, 8'd34}: color_data = 12'h000;
			{8'd106, 8'd35}: color_data = 12'h000;
			{8'd106, 8'd36}: color_data = 12'h000;
			{8'd106, 8'd37}: color_data = 12'h000;
			{8'd106, 8'd38}: color_data = 12'h980;
			{8'd106, 8'd39}: color_data = 12'hfd0;
			{8'd106, 8'd40}: color_data = 12'hfc0;
			{8'd106, 8'd41}: color_data = 12'hfc0;
			{8'd106, 8'd42}: color_data = 12'hfc0;
			{8'd106, 8'd43}: color_data = 12'hfc0;
			{8'd106, 8'd44}: color_data = 12'hfc0;
			{8'd106, 8'd45}: color_data = 12'hfc0;
			{8'd106, 8'd46}: color_data = 12'hfc0;
			{8'd106, 8'd47}: color_data = 12'hfc0;
			{8'd106, 8'd48}: color_data = 12'hfc0;
			{8'd106, 8'd49}: color_data = 12'hfd0;
			{8'd106, 8'd50}: color_data = 12'hfd0;
			{8'd106, 8'd51}: color_data = 12'hfd0;
			{8'd106, 8'd52}: color_data = 12'h870;
			{8'd106, 8'd53}: color_data = 12'h000;
			{8'd106, 8'd54}: color_data = 12'h000;
			{8'd106, 8'd55}: color_data = 12'h000;
			{8'd106, 8'd56}: color_data = 12'h000;
			{8'd106, 8'd57}: color_data = 12'h000;
			{8'd106, 8'd58}: color_data = 12'h000;
			{8'd106, 8'd59}: color_data = 12'h540;
			{8'd106, 8'd60}: color_data = 12'hfc0;
			{8'd106, 8'd61}: color_data = 12'hfd0;
			{8'd106, 8'd62}: color_data = 12'hfc0;
			{8'd106, 8'd63}: color_data = 12'hfc0;
			{8'd106, 8'd64}: color_data = 12'hfd0;
			{8'd106, 8'd65}: color_data = 12'h750;
			{8'd106, 8'd66}: color_data = 12'h000;
			{8'd106, 8'd67}: color_data = 12'h000;
			{8'd106, 8'd68}: color_data = 12'h000;
			{8'd106, 8'd69}: color_data = 12'h000;
			{8'd106, 8'd70}: color_data = 12'h000;
			{8'd106, 8'd71}: color_data = 12'h000;
			{8'd106, 8'd72}: color_data = 12'h000;
			{8'd106, 8'd100}: color_data = 12'he00;
			{8'd106, 8'd101}: color_data = 12'hf01;
			{8'd106, 8'd102}: color_data = 12'he00;
			{8'd106, 8'd103}: color_data = 12'he00;
			{8'd106, 8'd104}: color_data = 12'he00;
			{8'd106, 8'd105}: color_data = 12'he00;
			{8'd106, 8'd106}: color_data = 12'hc00;
			{8'd106, 8'd118}: color_data = 12'he00;
			{8'd106, 8'd119}: color_data = 12'he00;
			{8'd106, 8'd120}: color_data = 12'he00;
			{8'd106, 8'd121}: color_data = 12'he00;
			{8'd106, 8'd122}: color_data = 12'he00;
			{8'd106, 8'd123}: color_data = 12'he00;
			{8'd106, 8'd124}: color_data = 12'he00;
			{8'd106, 8'd125}: color_data = 12'he00;
			{8'd106, 8'd126}: color_data = 12'he00;
			{8'd106, 8'd127}: color_data = 12'he00;
			{8'd106, 8'd128}: color_data = 12'he00;
			{8'd106, 8'd129}: color_data = 12'he00;
			{8'd106, 8'd130}: color_data = 12'he00;
			{8'd106, 8'd131}: color_data = 12'hf01;
			{8'd106, 8'd132}: color_data = 12'he00;
			{8'd106, 8'd133}: color_data = 12'he01;
			{8'd106, 8'd138}: color_data = 12'he00;
			{8'd106, 8'd139}: color_data = 12'he00;
			{8'd106, 8'd140}: color_data = 12'he00;
			{8'd106, 8'd141}: color_data = 12'he00;
			{8'd106, 8'd142}: color_data = 12'he00;
			{8'd106, 8'd143}: color_data = 12'he01;
			{8'd106, 8'd144}: color_data = 12'he00;
			{8'd107, 8'd3}: color_data = 12'h000;
			{8'd107, 8'd4}: color_data = 12'h000;
			{8'd107, 8'd5}: color_data = 12'h131;
			{8'd107, 8'd6}: color_data = 12'h4b3;
			{8'd107, 8'd7}: color_data = 12'h4a3;
			{8'd107, 8'd8}: color_data = 12'h4a3;
			{8'd107, 8'd9}: color_data = 12'h4a3;
			{8'd107, 8'd10}: color_data = 12'h4a3;
			{8'd107, 8'd11}: color_data = 12'h4a3;
			{8'd107, 8'd12}: color_data = 12'h4b3;
			{8'd107, 8'd13}: color_data = 12'h4b3;
			{8'd107, 8'd14}: color_data = 12'h4b3;
			{8'd107, 8'd15}: color_data = 12'h4b3;
			{8'd107, 8'd16}: color_data = 12'h4a3;
			{8'd107, 8'd17}: color_data = 12'h4a3;
			{8'd107, 8'd18}: color_data = 12'h4a3;
			{8'd107, 8'd19}: color_data = 12'h4b3;
			{8'd107, 8'd20}: color_data = 12'h392;
			{8'd107, 8'd21}: color_data = 12'h392;
			{8'd107, 8'd22}: color_data = 12'h4a3;
			{8'd107, 8'd23}: color_data = 12'h4b3;
			{8'd107, 8'd24}: color_data = 12'h4b3;
			{8'd107, 8'd25}: color_data = 12'h4a3;
			{8'd107, 8'd26}: color_data = 12'h4a3;
			{8'd107, 8'd27}: color_data = 12'h4a3;
			{8'd107, 8'd28}: color_data = 12'h4b3;
			{8'd107, 8'd29}: color_data = 12'h3a3;
			{8'd107, 8'd30}: color_data = 12'h010;
			{8'd107, 8'd31}: color_data = 12'h000;
			{8'd107, 8'd32}: color_data = 12'h000;
			{8'd107, 8'd33}: color_data = 12'h000;
			{8'd107, 8'd34}: color_data = 12'h000;
			{8'd107, 8'd35}: color_data = 12'h000;
			{8'd107, 8'd36}: color_data = 12'h000;
			{8'd107, 8'd37}: color_data = 12'h000;
			{8'd107, 8'd38}: color_data = 12'h210;
			{8'd107, 8'd39}: color_data = 12'heb0;
			{8'd107, 8'd40}: color_data = 12'hfd0;
			{8'd107, 8'd41}: color_data = 12'hfc0;
			{8'd107, 8'd42}: color_data = 12'hfc0;
			{8'd107, 8'd43}: color_data = 12'hfc0;
			{8'd107, 8'd44}: color_data = 12'hfd0;
			{8'd107, 8'd45}: color_data = 12'hfd0;
			{8'd107, 8'd46}: color_data = 12'hfd0;
			{8'd107, 8'd47}: color_data = 12'hfd0;
			{8'd107, 8'd48}: color_data = 12'hfd0;
			{8'd107, 8'd49}: color_data = 12'hfc0;
			{8'd107, 8'd50}: color_data = 12'hdb0;
			{8'd107, 8'd51}: color_data = 12'ha80;
			{8'd107, 8'd52}: color_data = 12'h110;
			{8'd107, 8'd53}: color_data = 12'h000;
			{8'd107, 8'd54}: color_data = 12'h000;
			{8'd107, 8'd55}: color_data = 12'h000;
			{8'd107, 8'd56}: color_data = 12'h000;
			{8'd107, 8'd57}: color_data = 12'h000;
			{8'd107, 8'd58}: color_data = 12'h000;
			{8'd107, 8'd59}: color_data = 12'h000;
			{8'd107, 8'd60}: color_data = 12'h760;
			{8'd107, 8'd61}: color_data = 12'hfd0;
			{8'd107, 8'd62}: color_data = 12'hfd0;
			{8'd107, 8'd63}: color_data = 12'hfd0;
			{8'd107, 8'd64}: color_data = 12'heb0;
			{8'd107, 8'd65}: color_data = 12'h110;
			{8'd107, 8'd66}: color_data = 12'h000;
			{8'd107, 8'd67}: color_data = 12'h000;
			{8'd107, 8'd68}: color_data = 12'h000;
			{8'd107, 8'd69}: color_data = 12'h000;
			{8'd107, 8'd70}: color_data = 12'h000;
			{8'd107, 8'd71}: color_data = 12'h000;
			{8'd107, 8'd72}: color_data = 12'h000;
			{8'd107, 8'd100}: color_data = 12'he00;
			{8'd107, 8'd101}: color_data = 12'hf01;
			{8'd107, 8'd102}: color_data = 12'he00;
			{8'd107, 8'd103}: color_data = 12'he00;
			{8'd107, 8'd104}: color_data = 12'he00;
			{8'd107, 8'd105}: color_data = 12'he00;
			{8'd107, 8'd106}: color_data = 12'hc00;
			{8'd107, 8'd117}: color_data = 12'hd00;
			{8'd107, 8'd118}: color_data = 12'he00;
			{8'd107, 8'd119}: color_data = 12'he00;
			{8'd107, 8'd120}: color_data = 12'he00;
			{8'd107, 8'd121}: color_data = 12'he00;
			{8'd107, 8'd122}: color_data = 12'he00;
			{8'd107, 8'd123}: color_data = 12'he00;
			{8'd107, 8'd124}: color_data = 12'he00;
			{8'd107, 8'd125}: color_data = 12'he00;
			{8'd107, 8'd126}: color_data = 12'he00;
			{8'd107, 8'd127}: color_data = 12'he00;
			{8'd107, 8'd128}: color_data = 12'he00;
			{8'd107, 8'd129}: color_data = 12'he00;
			{8'd107, 8'd130}: color_data = 12'he00;
			{8'd107, 8'd131}: color_data = 12'he00;
			{8'd107, 8'd132}: color_data = 12'hf00;
			{8'd107, 8'd133}: color_data = 12'he00;
			{8'd107, 8'd138}: color_data = 12'he00;
			{8'd107, 8'd139}: color_data = 12'he00;
			{8'd107, 8'd140}: color_data = 12'he00;
			{8'd107, 8'd141}: color_data = 12'he00;
			{8'd107, 8'd142}: color_data = 12'he00;
			{8'd107, 8'd143}: color_data = 12'he01;
			{8'd107, 8'd144}: color_data = 12'he00;
			{8'd108, 8'd3}: color_data = 12'h000;
			{8'd108, 8'd4}: color_data = 12'h000;
			{8'd108, 8'd5}: color_data = 12'h020;
			{8'd108, 8'd6}: color_data = 12'h4a3;
			{8'd108, 8'd7}: color_data = 12'h4b3;
			{8'd108, 8'd8}: color_data = 12'h4a3;
			{8'd108, 8'd9}: color_data = 12'h4a3;
			{8'd108, 8'd10}: color_data = 12'h4a3;
			{8'd108, 8'd11}: color_data = 12'h4b3;
			{8'd108, 8'd12}: color_data = 12'h4a3;
			{8'd108, 8'd13}: color_data = 12'h392;
			{8'd108, 8'd14}: color_data = 12'h262;
			{8'd108, 8'd15}: color_data = 12'h251;
			{8'd108, 8'd16}: color_data = 12'h4a3;
			{8'd108, 8'd17}: color_data = 12'h4b3;
			{8'd108, 8'd18}: color_data = 12'h4a3;
			{8'd108, 8'd19}: color_data = 12'h4b3;
			{8'd108, 8'd20}: color_data = 12'h141;
			{8'd108, 8'd21}: color_data = 12'h000;
			{8'd108, 8'd22}: color_data = 12'h010;
			{8'd108, 8'd23}: color_data = 12'h120;
			{8'd108, 8'd24}: color_data = 12'h251;
			{8'd108, 8'd25}: color_data = 12'h4b3;
			{8'd108, 8'd26}: color_data = 12'h4a3;
			{8'd108, 8'd27}: color_data = 12'h4a3;
			{8'd108, 8'd28}: color_data = 12'h4b3;
			{8'd108, 8'd29}: color_data = 12'h4a3;
			{8'd108, 8'd30}: color_data = 12'h010;
			{8'd108, 8'd31}: color_data = 12'h000;
			{8'd108, 8'd32}: color_data = 12'h000;
			{8'd108, 8'd33}: color_data = 12'h000;
			{8'd108, 8'd34}: color_data = 12'h000;
			{8'd108, 8'd35}: color_data = 12'h000;
			{8'd108, 8'd36}: color_data = 12'h000;
			{8'd108, 8'd37}: color_data = 12'h000;
			{8'd108, 8'd38}: color_data = 12'h000;
			{8'd108, 8'd39}: color_data = 12'h760;
			{8'd108, 8'd40}: color_data = 12'hfd0;
			{8'd108, 8'd41}: color_data = 12'hfd0;
			{8'd108, 8'd42}: color_data = 12'hfd0;
			{8'd108, 8'd43}: color_data = 12'hfd0;
			{8'd108, 8'd44}: color_data = 12'hfc0;
			{8'd108, 8'd45}: color_data = 12'hda0;
			{8'd108, 8'd46}: color_data = 12'ha80;
			{8'd108, 8'd47}: color_data = 12'h760;
			{8'd108, 8'd48}: color_data = 12'h540;
			{8'd108, 8'd49}: color_data = 12'h220;
			{8'd108, 8'd50}: color_data = 12'h000;
			{8'd108, 8'd51}: color_data = 12'h000;
			{8'd108, 8'd52}: color_data = 12'h000;
			{8'd108, 8'd53}: color_data = 12'h000;
			{8'd108, 8'd54}: color_data = 12'h000;
			{8'd108, 8'd55}: color_data = 12'h000;
			{8'd108, 8'd56}: color_data = 12'h000;
			{8'd108, 8'd57}: color_data = 12'h000;
			{8'd108, 8'd58}: color_data = 12'h000;
			{8'd108, 8'd59}: color_data = 12'h000;
			{8'd108, 8'd60}: color_data = 12'h000;
			{8'd108, 8'd61}: color_data = 12'h970;
			{8'd108, 8'd62}: color_data = 12'hfd0;
			{8'd108, 8'd63}: color_data = 12'hfd0;
			{8'd108, 8'd64}: color_data = 12'h870;
			{8'd108, 8'd65}: color_data = 12'h000;
			{8'd108, 8'd66}: color_data = 12'h000;
			{8'd108, 8'd67}: color_data = 12'h000;
			{8'd108, 8'd68}: color_data = 12'h000;
			{8'd108, 8'd69}: color_data = 12'h000;
			{8'd108, 8'd70}: color_data = 12'h000;
			{8'd108, 8'd71}: color_data = 12'h000;
			{8'd108, 8'd73}: color_data = 12'h000;
			{8'd108, 8'd74}: color_data = 12'h000;
			{8'd108, 8'd100}: color_data = 12'he00;
			{8'd108, 8'd101}: color_data = 12'hf01;
			{8'd108, 8'd102}: color_data = 12'he00;
			{8'd108, 8'd103}: color_data = 12'he00;
			{8'd108, 8'd104}: color_data = 12'he00;
			{8'd108, 8'd105}: color_data = 12'he00;
			{8'd108, 8'd106}: color_data = 12'hc00;
			{8'd108, 8'd117}: color_data = 12'he00;
			{8'd108, 8'd118}: color_data = 12'he00;
			{8'd108, 8'd119}: color_data = 12'he00;
			{8'd108, 8'd120}: color_data = 12'he00;
			{8'd108, 8'd121}: color_data = 12'he00;
			{8'd108, 8'd122}: color_data = 12'he00;
			{8'd108, 8'd123}: color_data = 12'he00;
			{8'd108, 8'd124}: color_data = 12'he01;
			{8'd108, 8'd125}: color_data = 12'he01;
			{8'd108, 8'd126}: color_data = 12'he01;
			{8'd108, 8'd127}: color_data = 12'he01;
			{8'd108, 8'd128}: color_data = 12'he00;
			{8'd108, 8'd129}: color_data = 12'he00;
			{8'd108, 8'd130}: color_data = 12'he00;
			{8'd108, 8'd131}: color_data = 12'he00;
			{8'd108, 8'd132}: color_data = 12'he00;
			{8'd108, 8'd133}: color_data = 12'he00;
			{8'd108, 8'd138}: color_data = 12'he00;
			{8'd108, 8'd139}: color_data = 12'he00;
			{8'd108, 8'd140}: color_data = 12'he00;
			{8'd108, 8'd141}: color_data = 12'he00;
			{8'd108, 8'd142}: color_data = 12'he00;
			{8'd108, 8'd143}: color_data = 12'he01;
			{8'd108, 8'd144}: color_data = 12'he00;
			{8'd109, 8'd3}: color_data = 12'h000;
			{8'd109, 8'd4}: color_data = 12'h000;
			{8'd109, 8'd5}: color_data = 12'h000;
			{8'd109, 8'd6}: color_data = 12'h393;
			{8'd109, 8'd7}: color_data = 12'h4b3;
			{8'd109, 8'd8}: color_data = 12'h4a3;
			{8'd109, 8'd9}: color_data = 12'h4a3;
			{8'd109, 8'd10}: color_data = 12'h4b3;
			{8'd109, 8'd11}: color_data = 12'h392;
			{8'd109, 8'd12}: color_data = 12'h020;
			{8'd109, 8'd13}: color_data = 12'h000;
			{8'd109, 8'd14}: color_data = 12'h000;
			{8'd109, 8'd15}: color_data = 12'h010;
			{8'd109, 8'd16}: color_data = 12'h4a3;
			{8'd109, 8'd17}: color_data = 12'h4b3;
			{8'd109, 8'd18}: color_data = 12'h4a3;
			{8'd109, 8'd19}: color_data = 12'h4b3;
			{8'd109, 8'd20}: color_data = 12'h261;
			{8'd109, 8'd21}: color_data = 12'h000;
			{8'd109, 8'd22}: color_data = 12'h000;
			{8'd109, 8'd23}: color_data = 12'h000;
			{8'd109, 8'd24}: color_data = 12'h141;
			{8'd109, 8'd25}: color_data = 12'h4b3;
			{8'd109, 8'd26}: color_data = 12'h4a3;
			{8'd109, 8'd27}: color_data = 12'h4a3;
			{8'd109, 8'd28}: color_data = 12'h4b3;
			{8'd109, 8'd29}: color_data = 12'h4a3;
			{8'd109, 8'd30}: color_data = 12'h010;
			{8'd109, 8'd31}: color_data = 12'h000;
			{8'd109, 8'd32}: color_data = 12'h000;
			{8'd109, 8'd33}: color_data = 12'h000;
			{8'd109, 8'd34}: color_data = 12'h000;
			{8'd109, 8'd35}: color_data = 12'h000;
			{8'd109, 8'd36}: color_data = 12'h000;
			{8'd109, 8'd37}: color_data = 12'h000;
			{8'd109, 8'd38}: color_data = 12'h000;
			{8'd109, 8'd39}: color_data = 12'h000;
			{8'd109, 8'd40}: color_data = 12'ha80;
			{8'd109, 8'd41}: color_data = 12'ha80;
			{8'd109, 8'd42}: color_data = 12'h760;
			{8'd109, 8'd43}: color_data = 12'h430;
			{8'd109, 8'd44}: color_data = 12'h210;
			{8'd109, 8'd45}: color_data = 12'h000;
			{8'd109, 8'd46}: color_data = 12'h000;
			{8'd109, 8'd47}: color_data = 12'h000;
			{8'd109, 8'd48}: color_data = 12'h000;
			{8'd109, 8'd49}: color_data = 12'h000;
			{8'd109, 8'd50}: color_data = 12'h000;
			{8'd109, 8'd51}: color_data = 12'h000;
			{8'd109, 8'd52}: color_data = 12'h000;
			{8'd109, 8'd53}: color_data = 12'h000;
			{8'd109, 8'd54}: color_data = 12'h000;
			{8'd109, 8'd55}: color_data = 12'h000;
			{8'd109, 8'd56}: color_data = 12'h000;
			{8'd109, 8'd57}: color_data = 12'h000;
			{8'd109, 8'd58}: color_data = 12'h000;
			{8'd109, 8'd59}: color_data = 12'h000;
			{8'd109, 8'd60}: color_data = 12'h000;
			{8'd109, 8'd61}: color_data = 12'h000;
			{8'd109, 8'd62}: color_data = 12'hb90;
			{8'd109, 8'd63}: color_data = 12'hfd0;
			{8'd109, 8'd64}: color_data = 12'h220;
			{8'd109, 8'd65}: color_data = 12'h000;
			{8'd109, 8'd66}: color_data = 12'h000;
			{8'd109, 8'd67}: color_data = 12'h000;
			{8'd109, 8'd68}: color_data = 12'h000;
			{8'd109, 8'd69}: color_data = 12'h000;
			{8'd109, 8'd70}: color_data = 12'h000;
			{8'd109, 8'd71}: color_data = 12'h000;
			{8'd109, 8'd72}: color_data = 12'h000;
			{8'd109, 8'd73}: color_data = 12'h000;
			{8'd109, 8'd74}: color_data = 12'h000;
			{8'd109, 8'd75}: color_data = 12'h000;
			{8'd109, 8'd100}: color_data = 12'he00;
			{8'd109, 8'd101}: color_data = 12'hf01;
			{8'd109, 8'd102}: color_data = 12'he00;
			{8'd109, 8'd103}: color_data = 12'he00;
			{8'd109, 8'd104}: color_data = 12'he00;
			{8'd109, 8'd105}: color_data = 12'he00;
			{8'd109, 8'd106}: color_data = 12'hc00;
			{8'd109, 8'd117}: color_data = 12'he00;
			{8'd109, 8'd118}: color_data = 12'he01;
			{8'd109, 8'd119}: color_data = 12'he00;
			{8'd109, 8'd120}: color_data = 12'he00;
			{8'd109, 8'd121}: color_data = 12'he00;
			{8'd109, 8'd122}: color_data = 12'he00;
			{8'd109, 8'd123}: color_data = 12'he00;
			{8'd109, 8'd124}: color_data = 12'he00;
			{8'd109, 8'd125}: color_data = 12'he00;
			{8'd109, 8'd126}: color_data = 12'he00;
			{8'd109, 8'd127}: color_data = 12'he00;
			{8'd109, 8'd128}: color_data = 12'he00;
			{8'd109, 8'd129}: color_data = 12'he00;
			{8'd109, 8'd130}: color_data = 12'he00;
			{8'd109, 8'd131}: color_data = 12'he00;
			{8'd109, 8'd132}: color_data = 12'he00;
			{8'd109, 8'd133}: color_data = 12'he00;
			{8'd109, 8'd134}: color_data = 12'hd00;
			{8'd109, 8'd138}: color_data = 12'he00;
			{8'd109, 8'd139}: color_data = 12'he00;
			{8'd109, 8'd140}: color_data = 12'he00;
			{8'd109, 8'd141}: color_data = 12'he00;
			{8'd109, 8'd142}: color_data = 12'he00;
			{8'd109, 8'd143}: color_data = 12'he01;
			{8'd109, 8'd144}: color_data = 12'he00;
			{8'd110, 8'd3}: color_data = 12'h000;
			{8'd110, 8'd4}: color_data = 12'h000;
			{8'd110, 8'd5}: color_data = 12'h000;
			{8'd110, 8'd6}: color_data = 12'h382;
			{8'd110, 8'd7}: color_data = 12'h4b3;
			{8'd110, 8'd8}: color_data = 12'h4a3;
			{8'd110, 8'd9}: color_data = 12'h4a3;
			{8'd110, 8'd10}: color_data = 12'h4b3;
			{8'd110, 8'd11}: color_data = 12'h3a3;
			{8'd110, 8'd12}: color_data = 12'h010;
			{8'd110, 8'd13}: color_data = 12'h000;
			{8'd110, 8'd14}: color_data = 12'h000;
			{8'd110, 8'd15}: color_data = 12'h010;
			{8'd110, 8'd16}: color_data = 12'h4a3;
			{8'd110, 8'd17}: color_data = 12'h4b3;
			{8'd110, 8'd18}: color_data = 12'h4a3;
			{8'd110, 8'd19}: color_data = 12'h4b3;
			{8'd110, 8'd20}: color_data = 12'h372;
			{8'd110, 8'd21}: color_data = 12'h000;
			{8'd110, 8'd22}: color_data = 12'h000;
			{8'd110, 8'd23}: color_data = 12'h000;
			{8'd110, 8'd24}: color_data = 12'h251;
			{8'd110, 8'd25}: color_data = 12'h4b3;
			{8'd110, 8'd26}: color_data = 12'h4a3;
			{8'd110, 8'd27}: color_data = 12'h4a3;
			{8'd110, 8'd28}: color_data = 12'h4b3;
			{8'd110, 8'd29}: color_data = 12'h4a3;
			{8'd110, 8'd30}: color_data = 12'h010;
			{8'd110, 8'd31}: color_data = 12'h000;
			{8'd110, 8'd32}: color_data = 12'h000;
			{8'd110, 8'd33}: color_data = 12'h000;
			{8'd110, 8'd34}: color_data = 12'h000;
			{8'd110, 8'd35}: color_data = 12'h000;
			{8'd110, 8'd36}: color_data = 12'h000;
			{8'd110, 8'd37}: color_data = 12'h000;
			{8'd110, 8'd38}: color_data = 12'h000;
			{8'd110, 8'd39}: color_data = 12'h000;
			{8'd110, 8'd40}: color_data = 12'h000;
			{8'd110, 8'd41}: color_data = 12'h000;
			{8'd110, 8'd42}: color_data = 12'h000;
			{8'd110, 8'd43}: color_data = 12'h000;
			{8'd110, 8'd44}: color_data = 12'h000;
			{8'd110, 8'd45}: color_data = 12'h000;
			{8'd110, 8'd46}: color_data = 12'h000;
			{8'd110, 8'd47}: color_data = 12'h000;
			{8'd110, 8'd48}: color_data = 12'h000;
			{8'd110, 8'd49}: color_data = 12'h000;
			{8'd110, 8'd50}: color_data = 12'h000;
			{8'd110, 8'd51}: color_data = 12'h000;
			{8'd110, 8'd52}: color_data = 12'h000;
			{8'd110, 8'd53}: color_data = 12'h000;
			{8'd110, 8'd54}: color_data = 12'h000;
			{8'd110, 8'd55}: color_data = 12'h000;
			{8'd110, 8'd56}: color_data = 12'h000;
			{8'd110, 8'd57}: color_data = 12'h000;
			{8'd110, 8'd58}: color_data = 12'h000;
			{8'd110, 8'd59}: color_data = 12'h000;
			{8'd110, 8'd60}: color_data = 12'h000;
			{8'd110, 8'd61}: color_data = 12'h000;
			{8'd110, 8'd62}: color_data = 12'h210;
			{8'd110, 8'd63}: color_data = 12'h750;
			{8'd110, 8'd64}: color_data = 12'h000;
			{8'd110, 8'd65}: color_data = 12'h000;
			{8'd110, 8'd66}: color_data = 12'h000;
			{8'd110, 8'd67}: color_data = 12'h000;
			{8'd110, 8'd68}: color_data = 12'h000;
			{8'd110, 8'd69}: color_data = 12'h000;
			{8'd110, 8'd70}: color_data = 12'h000;
			{8'd110, 8'd71}: color_data = 12'h000;
			{8'd110, 8'd72}: color_data = 12'h000;
			{8'd110, 8'd73}: color_data = 12'h000;
			{8'd110, 8'd74}: color_data = 12'h000;
			{8'd110, 8'd75}: color_data = 12'h000;
			{8'd110, 8'd100}: color_data = 12'he00;
			{8'd110, 8'd101}: color_data = 12'hf01;
			{8'd110, 8'd102}: color_data = 12'he00;
			{8'd110, 8'd103}: color_data = 12'he00;
			{8'd110, 8'd104}: color_data = 12'he00;
			{8'd110, 8'd105}: color_data = 12'he00;
			{8'd110, 8'd106}: color_data = 12'hc00;
			{8'd110, 8'd117}: color_data = 12'he00;
			{8'd110, 8'd118}: color_data = 12'he01;
			{8'd110, 8'd119}: color_data = 12'he00;
			{8'd110, 8'd120}: color_data = 12'he00;
			{8'd110, 8'd121}: color_data = 12'he00;
			{8'd110, 8'd122}: color_data = 12'he00;
			{8'd110, 8'd123}: color_data = 12'hf00;
			{8'd110, 8'd128}: color_data = 12'he00;
			{8'd110, 8'd129}: color_data = 12'he00;
			{8'd110, 8'd130}: color_data = 12'he00;
			{8'd110, 8'd131}: color_data = 12'he00;
			{8'd110, 8'd132}: color_data = 12'he00;
			{8'd110, 8'd133}: color_data = 12'he00;
			{8'd110, 8'd134}: color_data = 12'hf00;
			{8'd110, 8'd138}: color_data = 12'he00;
			{8'd110, 8'd139}: color_data = 12'he00;
			{8'd110, 8'd140}: color_data = 12'he00;
			{8'd110, 8'd141}: color_data = 12'he00;
			{8'd110, 8'd142}: color_data = 12'he00;
			{8'd110, 8'd143}: color_data = 12'he01;
			{8'd110, 8'd144}: color_data = 12'he00;
			{8'd111, 8'd3}: color_data = 12'h000;
			{8'd111, 8'd4}: color_data = 12'h000;
			{8'd111, 8'd5}: color_data = 12'h000;
			{8'd111, 8'd6}: color_data = 12'h262;
			{8'd111, 8'd7}: color_data = 12'h4b3;
			{8'd111, 8'd8}: color_data = 12'h4a3;
			{8'd111, 8'd9}: color_data = 12'h4a3;
			{8'd111, 8'd10}: color_data = 12'h4a3;
			{8'd111, 8'd11}: color_data = 12'h4b3;
			{8'd111, 8'd12}: color_data = 12'h131;
			{8'd111, 8'd13}: color_data = 12'h000;
			{8'd111, 8'd14}: color_data = 12'h000;
			{8'd111, 8'd15}: color_data = 12'h010;
			{8'd111, 8'd16}: color_data = 12'h4a3;
			{8'd111, 8'd17}: color_data = 12'h4b3;
			{8'd111, 8'd18}: color_data = 12'h4a3;
			{8'd111, 8'd19}: color_data = 12'h4b3;
			{8'd111, 8'd20}: color_data = 12'h392;
			{8'd111, 8'd21}: color_data = 12'h000;
			{8'd111, 8'd22}: color_data = 12'h000;
			{8'd111, 8'd23}: color_data = 12'h000;
			{8'd111, 8'd24}: color_data = 12'h272;
			{8'd111, 8'd25}: color_data = 12'h4b3;
			{8'd111, 8'd26}: color_data = 12'h4a3;
			{8'd111, 8'd27}: color_data = 12'h4a3;
			{8'd111, 8'd28}: color_data = 12'h4b3;
			{8'd111, 8'd29}: color_data = 12'h4a3;
			{8'd111, 8'd30}: color_data = 12'h020;
			{8'd111, 8'd31}: color_data = 12'h000;
			{8'd111, 8'd32}: color_data = 12'h000;
			{8'd111, 8'd33}: color_data = 12'h000;
			{8'd111, 8'd34}: color_data = 12'h000;
			{8'd111, 8'd35}: color_data = 12'h000;
			{8'd111, 8'd36}: color_data = 12'h000;
			{8'd111, 8'd37}: color_data = 12'h000;
			{8'd111, 8'd38}: color_data = 12'h000;
			{8'd111, 8'd39}: color_data = 12'h000;
			{8'd111, 8'd40}: color_data = 12'h000;
			{8'd111, 8'd41}: color_data = 12'h000;
			{8'd111, 8'd42}: color_data = 12'h000;
			{8'd111, 8'd43}: color_data = 12'h000;
			{8'd111, 8'd44}: color_data = 12'h000;
			{8'd111, 8'd45}: color_data = 12'h000;
			{8'd111, 8'd46}: color_data = 12'h000;
			{8'd111, 8'd47}: color_data = 12'h000;
			{8'd111, 8'd48}: color_data = 12'h000;
			{8'd111, 8'd49}: color_data = 12'h000;
			{8'd111, 8'd50}: color_data = 12'h000;
			{8'd111, 8'd51}: color_data = 12'h000;
			{8'd111, 8'd52}: color_data = 12'h000;
			{8'd111, 8'd53}: color_data = 12'h000;
			{8'd111, 8'd54}: color_data = 12'h000;
			{8'd111, 8'd55}: color_data = 12'h000;
			{8'd111, 8'd56}: color_data = 12'h000;
			{8'd111, 8'd57}: color_data = 12'h000;
			{8'd111, 8'd58}: color_data = 12'h000;
			{8'd111, 8'd59}: color_data = 12'h000;
			{8'd111, 8'd60}: color_data = 12'h000;
			{8'd111, 8'd61}: color_data = 12'h000;
			{8'd111, 8'd62}: color_data = 12'h000;
			{8'd111, 8'd63}: color_data = 12'h000;
			{8'd111, 8'd64}: color_data = 12'h000;
			{8'd111, 8'd65}: color_data = 12'h000;
			{8'd111, 8'd66}: color_data = 12'h011;
			{8'd111, 8'd67}: color_data = 12'h011;
			{8'd111, 8'd68}: color_data = 12'h000;
			{8'd111, 8'd69}: color_data = 12'h000;
			{8'd111, 8'd70}: color_data = 12'h000;
			{8'd111, 8'd71}: color_data = 12'h000;
			{8'd111, 8'd72}: color_data = 12'h000;
			{8'd111, 8'd73}: color_data = 12'h000;
			{8'd111, 8'd74}: color_data = 12'h000;
			{8'd111, 8'd75}: color_data = 12'h000;
			{8'd111, 8'd100}: color_data = 12'he00;
			{8'd111, 8'd101}: color_data = 12'hf01;
			{8'd111, 8'd102}: color_data = 12'he00;
			{8'd111, 8'd103}: color_data = 12'he00;
			{8'd111, 8'd104}: color_data = 12'he00;
			{8'd111, 8'd105}: color_data = 12'he00;
			{8'd111, 8'd106}: color_data = 12'hc00;
			{8'd111, 8'd117}: color_data = 12'he00;
			{8'd111, 8'd118}: color_data = 12'he00;
			{8'd111, 8'd119}: color_data = 12'he00;
			{8'd111, 8'd120}: color_data = 12'he00;
			{8'd111, 8'd121}: color_data = 12'he00;
			{8'd111, 8'd122}: color_data = 12'he01;
			{8'd111, 8'd129}: color_data = 12'he00;
			{8'd111, 8'd130}: color_data = 12'he01;
			{8'd111, 8'd131}: color_data = 12'he00;
			{8'd111, 8'd132}: color_data = 12'he00;
			{8'd111, 8'd133}: color_data = 12'he00;
			{8'd111, 8'd138}: color_data = 12'he00;
			{8'd111, 8'd139}: color_data = 12'he00;
			{8'd111, 8'd140}: color_data = 12'he00;
			{8'd111, 8'd141}: color_data = 12'he00;
			{8'd111, 8'd142}: color_data = 12'he00;
			{8'd111, 8'd143}: color_data = 12'he01;
			{8'd111, 8'd144}: color_data = 12'he00;
			{8'd112, 8'd4}: color_data = 12'h000;
			{8'd112, 8'd5}: color_data = 12'h000;
			{8'd112, 8'd6}: color_data = 12'h141;
			{8'd112, 8'd7}: color_data = 12'h4b3;
			{8'd112, 8'd8}: color_data = 12'h4a3;
			{8'd112, 8'd9}: color_data = 12'h4a3;
			{8'd112, 8'd10}: color_data = 12'h4a3;
			{8'd112, 8'd11}: color_data = 12'h4b3;
			{8'd112, 8'd12}: color_data = 12'h272;
			{8'd112, 8'd13}: color_data = 12'h000;
			{8'd112, 8'd14}: color_data = 12'h000;
			{8'd112, 8'd15}: color_data = 12'h010;
			{8'd112, 8'd16}: color_data = 12'h4a3;
			{8'd112, 8'd17}: color_data = 12'h4b3;
			{8'd112, 8'd18}: color_data = 12'h4a3;
			{8'd112, 8'd19}: color_data = 12'h4b3;
			{8'd112, 8'd20}: color_data = 12'h4a3;
			{8'd112, 8'd21}: color_data = 12'h010;
			{8'd112, 8'd22}: color_data = 12'h000;
			{8'd112, 8'd23}: color_data = 12'h000;
			{8'd112, 8'd24}: color_data = 12'h382;
			{8'd112, 8'd25}: color_data = 12'h4b3;
			{8'd112, 8'd26}: color_data = 12'h4a3;
			{8'd112, 8'd27}: color_data = 12'h4a3;
			{8'd112, 8'd28}: color_data = 12'h4b3;
			{8'd112, 8'd29}: color_data = 12'h4b3;
			{8'd112, 8'd30}: color_data = 12'h020;
			{8'd112, 8'd31}: color_data = 12'h000;
			{8'd112, 8'd32}: color_data = 12'h000;
			{8'd112, 8'd33}: color_data = 12'h000;
			{8'd112, 8'd34}: color_data = 12'h000;
			{8'd112, 8'd35}: color_data = 12'h000;
			{8'd112, 8'd36}: color_data = 12'h000;
			{8'd112, 8'd37}: color_data = 12'h000;
			{8'd112, 8'd38}: color_data = 12'h000;
			{8'd112, 8'd39}: color_data = 12'h001;
			{8'd112, 8'd40}: color_data = 12'h011;
			{8'd112, 8'd41}: color_data = 12'h011;
			{8'd112, 8'd42}: color_data = 12'h012;
			{8'd112, 8'd43}: color_data = 12'h012;
			{8'd112, 8'd44}: color_data = 12'h023;
			{8'd112, 8'd45}: color_data = 12'h023;
			{8'd112, 8'd46}: color_data = 12'h023;
			{8'd112, 8'd47}: color_data = 12'h034;
			{8'd112, 8'd48}: color_data = 12'h034;
			{8'd112, 8'd49}: color_data = 12'h035;
			{8'd112, 8'd50}: color_data = 12'h045;
			{8'd112, 8'd51}: color_data = 12'h046;
			{8'd112, 8'd52}: color_data = 12'h046;
			{8'd112, 8'd53}: color_data = 12'h057;
			{8'd112, 8'd54}: color_data = 12'h057;
			{8'd112, 8'd55}: color_data = 12'h058;
			{8'd112, 8'd56}: color_data = 12'h068;
			{8'd112, 8'd57}: color_data = 12'h069;
			{8'd112, 8'd58}: color_data = 12'h069;
			{8'd112, 8'd59}: color_data = 12'h07a;
			{8'd112, 8'd60}: color_data = 12'h07a;
			{8'd112, 8'd61}: color_data = 12'h023;
			{8'd112, 8'd62}: color_data = 12'h000;
			{8'd112, 8'd63}: color_data = 12'h000;
			{8'd112, 8'd64}: color_data = 12'h000;
			{8'd112, 8'd65}: color_data = 12'h034;
			{8'd112, 8'd66}: color_data = 12'h09d;
			{8'd112, 8'd67}: color_data = 12'h09d;
			{8'd112, 8'd68}: color_data = 12'h023;
			{8'd112, 8'd69}: color_data = 12'h000;
			{8'd112, 8'd70}: color_data = 12'h000;
			{8'd112, 8'd71}: color_data = 12'h000;
			{8'd112, 8'd72}: color_data = 12'h000;
			{8'd112, 8'd73}: color_data = 12'h000;
			{8'd112, 8'd74}: color_data = 12'h000;
			{8'd112, 8'd75}: color_data = 12'h000;
			{8'd112, 8'd100}: color_data = 12'he00;
			{8'd112, 8'd101}: color_data = 12'hf01;
			{8'd112, 8'd102}: color_data = 12'he00;
			{8'd112, 8'd103}: color_data = 12'he00;
			{8'd112, 8'd104}: color_data = 12'he00;
			{8'd112, 8'd105}: color_data = 12'he00;
			{8'd112, 8'd106}: color_data = 12'hc00;
			{8'd112, 8'd117}: color_data = 12'he00;
			{8'd112, 8'd118}: color_data = 12'he00;
			{8'd112, 8'd119}: color_data = 12'he00;
			{8'd112, 8'd120}: color_data = 12'he00;
			{8'd112, 8'd121}: color_data = 12'he00;
			{8'd112, 8'd122}: color_data = 12'he00;
			{8'd112, 8'd129}: color_data = 12'he00;
			{8'd112, 8'd130}: color_data = 12'he01;
			{8'd112, 8'd131}: color_data = 12'he00;
			{8'd112, 8'd132}: color_data = 12'he01;
			{8'd112, 8'd133}: color_data = 12'he00;
			{8'd112, 8'd138}: color_data = 12'he00;
			{8'd112, 8'd139}: color_data = 12'he00;
			{8'd112, 8'd140}: color_data = 12'he00;
			{8'd112, 8'd141}: color_data = 12'he00;
			{8'd112, 8'd142}: color_data = 12'he00;
			{8'd112, 8'd143}: color_data = 12'he01;
			{8'd112, 8'd144}: color_data = 12'he00;
			{8'd113, 8'd4}: color_data = 12'h000;
			{8'd113, 8'd5}: color_data = 12'h000;
			{8'd113, 8'd6}: color_data = 12'h130;
			{8'd113, 8'd7}: color_data = 12'h4b3;
			{8'd113, 8'd8}: color_data = 12'h4a3;
			{8'd113, 8'd9}: color_data = 12'h4a3;
			{8'd113, 8'd10}: color_data = 12'h4a3;
			{8'd113, 8'd11}: color_data = 12'h4b3;
			{8'd113, 8'd12}: color_data = 12'h392;
			{8'd113, 8'd13}: color_data = 12'h000;
			{8'd113, 8'd14}: color_data = 12'h000;
			{8'd113, 8'd15}: color_data = 12'h010;
			{8'd113, 8'd16}: color_data = 12'h3a3;
			{8'd113, 8'd17}: color_data = 12'h4b3;
			{8'd113, 8'd18}: color_data = 12'h4a3;
			{8'd113, 8'd19}: color_data = 12'h4b3;
			{8'd113, 8'd20}: color_data = 12'h4a3;
			{8'd113, 8'd21}: color_data = 12'h020;
			{8'd113, 8'd22}: color_data = 12'h000;
			{8'd113, 8'd23}: color_data = 12'h000;
			{8'd113, 8'd24}: color_data = 12'h393;
			{8'd113, 8'd25}: color_data = 12'h4b3;
			{8'd113, 8'd26}: color_data = 12'h4a3;
			{8'd113, 8'd27}: color_data = 12'h4a3;
			{8'd113, 8'd28}: color_data = 12'h4a3;
			{8'd113, 8'd29}: color_data = 12'h4b3;
			{8'd113, 8'd30}: color_data = 12'h120;
			{8'd113, 8'd31}: color_data = 12'h000;
			{8'd113, 8'd32}: color_data = 12'h000;
			{8'd113, 8'd33}: color_data = 12'h000;
			{8'd113, 8'd34}: color_data = 12'h069;
			{8'd113, 8'd35}: color_data = 12'h08b;
			{8'd113, 8'd36}: color_data = 12'h08b;
			{8'd113, 8'd37}: color_data = 12'h08b;
			{8'd113, 8'd38}: color_data = 12'h08c;
			{8'd113, 8'd39}: color_data = 12'h08c;
			{8'd113, 8'd40}: color_data = 12'h09c;
			{8'd113, 8'd41}: color_data = 12'h09c;
			{8'd113, 8'd42}: color_data = 12'h09d;
			{8'd113, 8'd43}: color_data = 12'h09d;
			{8'd113, 8'd44}: color_data = 12'h09d;
			{8'd113, 8'd45}: color_data = 12'h09d;
			{8'd113, 8'd46}: color_data = 12'h09d;
			{8'd113, 8'd47}: color_data = 12'h09d;
			{8'd113, 8'd48}: color_data = 12'h0ae;
			{8'd113, 8'd49}: color_data = 12'h0ae;
			{8'd113, 8'd50}: color_data = 12'h0ae;
			{8'd113, 8'd51}: color_data = 12'h0ae;
			{8'd113, 8'd52}: color_data = 12'h0ae;
			{8'd113, 8'd53}: color_data = 12'h0ae;
			{8'd113, 8'd54}: color_data = 12'h0ae;
			{8'd113, 8'd55}: color_data = 12'h0ae;
			{8'd113, 8'd56}: color_data = 12'h0ae;
			{8'd113, 8'd57}: color_data = 12'h0ae;
			{8'd113, 8'd58}: color_data = 12'h0ae;
			{8'd113, 8'd59}: color_data = 12'h0ae;
			{8'd113, 8'd60}: color_data = 12'h0ae;
			{8'd113, 8'd61}: color_data = 12'h08c;
			{8'd113, 8'd62}: color_data = 12'h023;
			{8'd113, 8'd63}: color_data = 12'h001;
			{8'd113, 8'd64}: color_data = 12'h022;
			{8'd113, 8'd65}: color_data = 12'h08b;
			{8'd113, 8'd66}: color_data = 12'h0ae;
			{8'd113, 8'd67}: color_data = 12'h09d;
			{8'd113, 8'd68}: color_data = 12'h023;
			{8'd113, 8'd69}: color_data = 12'h000;
			{8'd113, 8'd70}: color_data = 12'h000;
			{8'd113, 8'd71}: color_data = 12'h000;
			{8'd113, 8'd72}: color_data = 12'h000;
			{8'd113, 8'd73}: color_data = 12'h000;
			{8'd113, 8'd74}: color_data = 12'h000;
			{8'd113, 8'd75}: color_data = 12'h000;
			{8'd113, 8'd100}: color_data = 12'he00;
			{8'd113, 8'd101}: color_data = 12'hf01;
			{8'd113, 8'd102}: color_data = 12'he00;
			{8'd113, 8'd103}: color_data = 12'he00;
			{8'd113, 8'd104}: color_data = 12'he00;
			{8'd113, 8'd105}: color_data = 12'he00;
			{8'd113, 8'd106}: color_data = 12'hc00;
			{8'd113, 8'd118}: color_data = 12'he00;
			{8'd113, 8'd119}: color_data = 12'he00;
			{8'd113, 8'd120}: color_data = 12'he00;
			{8'd113, 8'd121}: color_data = 12'he00;
			{8'd113, 8'd122}: color_data = 12'he00;
			{8'd113, 8'd128}: color_data = 12'he00;
			{8'd113, 8'd129}: color_data = 12'he00;
			{8'd113, 8'd130}: color_data = 12'he00;
			{8'd113, 8'd131}: color_data = 12'he00;
			{8'd113, 8'd132}: color_data = 12'he00;
			{8'd113, 8'd133}: color_data = 12'hd00;
			{8'd113, 8'd138}: color_data = 12'he00;
			{8'd113, 8'd139}: color_data = 12'he00;
			{8'd113, 8'd140}: color_data = 12'he00;
			{8'd113, 8'd141}: color_data = 12'he00;
			{8'd113, 8'd142}: color_data = 12'he00;
			{8'd113, 8'd143}: color_data = 12'he01;
			{8'd113, 8'd144}: color_data = 12'he00;
			{8'd114, 8'd4}: color_data = 12'h000;
			{8'd114, 8'd5}: color_data = 12'h000;
			{8'd114, 8'd6}: color_data = 12'h010;
			{8'd114, 8'd7}: color_data = 12'h4a3;
			{8'd114, 8'd8}: color_data = 12'h4b3;
			{8'd114, 8'd9}: color_data = 12'h4a3;
			{8'd114, 8'd10}: color_data = 12'h4a3;
			{8'd114, 8'd11}: color_data = 12'h4b3;
			{8'd114, 8'd12}: color_data = 12'h4b3;
			{8'd114, 8'd13}: color_data = 12'h120;
			{8'd114, 8'd14}: color_data = 12'h000;
			{8'd114, 8'd15}: color_data = 12'h010;
			{8'd114, 8'd16}: color_data = 12'h4a3;
			{8'd114, 8'd17}: color_data = 12'h4b3;
			{8'd114, 8'd18}: color_data = 12'h4b3;
			{8'd114, 8'd19}: color_data = 12'h4b3;
			{8'd114, 8'd20}: color_data = 12'h4b3;
			{8'd114, 8'd21}: color_data = 12'h141;
			{8'd114, 8'd22}: color_data = 12'h000;
			{8'd114, 8'd23}: color_data = 12'h010;
			{8'd114, 8'd24}: color_data = 12'h4a3;
			{8'd114, 8'd25}: color_data = 12'h4b3;
			{8'd114, 8'd26}: color_data = 12'h4a3;
			{8'd114, 8'd27}: color_data = 12'h4a3;
			{8'd114, 8'd28}: color_data = 12'h4a3;
			{8'd114, 8'd29}: color_data = 12'h4b3;
			{8'd114, 8'd30}: color_data = 12'h130;
			{8'd114, 8'd31}: color_data = 12'h000;
			{8'd114, 8'd32}: color_data = 12'h000;
			{8'd114, 8'd33}: color_data = 12'h000;
			{8'd114, 8'd34}: color_data = 12'h08b;
			{8'd114, 8'd35}: color_data = 12'h0ae;
			{8'd114, 8'd36}: color_data = 12'h09d;
			{8'd114, 8'd37}: color_data = 12'h09d;
			{8'd114, 8'd38}: color_data = 12'h09d;
			{8'd114, 8'd39}: color_data = 12'h09d;
			{8'd114, 8'd40}: color_data = 12'h09d;
			{8'd114, 8'd41}: color_data = 12'h09d;
			{8'd114, 8'd42}: color_data = 12'h09d;
			{8'd114, 8'd43}: color_data = 12'h09d;
			{8'd114, 8'd44}: color_data = 12'h09d;
			{8'd114, 8'd45}: color_data = 12'h09d;
			{8'd114, 8'd46}: color_data = 12'h09d;
			{8'd114, 8'd47}: color_data = 12'h09d;
			{8'd114, 8'd48}: color_data = 12'h09d;
			{8'd114, 8'd49}: color_data = 12'h09d;
			{8'd114, 8'd50}: color_data = 12'h09d;
			{8'd114, 8'd51}: color_data = 12'h09d;
			{8'd114, 8'd52}: color_data = 12'h09d;
			{8'd114, 8'd53}: color_data = 12'h09d;
			{8'd114, 8'd54}: color_data = 12'h09d;
			{8'd114, 8'd55}: color_data = 12'h09d;
			{8'd114, 8'd56}: color_data = 12'h09d;
			{8'd114, 8'd57}: color_data = 12'h09d;
			{8'd114, 8'd58}: color_data = 12'h09d;
			{8'd114, 8'd59}: color_data = 12'h09d;
			{8'd114, 8'd60}: color_data = 12'h09d;
			{8'd114, 8'd61}: color_data = 12'h09d;
			{8'd114, 8'd62}: color_data = 12'h09d;
			{8'd114, 8'd63}: color_data = 12'h09c;
			{8'd114, 8'd64}: color_data = 12'h09d;
			{8'd114, 8'd65}: color_data = 12'h09d;
			{8'd114, 8'd66}: color_data = 12'h09d;
			{8'd114, 8'd67}: color_data = 12'h09d;
			{8'd114, 8'd68}: color_data = 12'h012;
			{8'd114, 8'd69}: color_data = 12'h000;
			{8'd114, 8'd70}: color_data = 12'h000;
			{8'd114, 8'd71}: color_data = 12'h000;
			{8'd114, 8'd72}: color_data = 12'h000;
			{8'd114, 8'd73}: color_data = 12'h000;
			{8'd114, 8'd74}: color_data = 12'h000;
			{8'd114, 8'd75}: color_data = 12'h000;
			{8'd114, 8'd100}: color_data = 12'he00;
			{8'd114, 8'd101}: color_data = 12'hf01;
			{8'd114, 8'd102}: color_data = 12'he00;
			{8'd114, 8'd103}: color_data = 12'he00;
			{8'd114, 8'd104}: color_data = 12'he00;
			{8'd114, 8'd105}: color_data = 12'he00;
			{8'd114, 8'd106}: color_data = 12'hc00;
			{8'd114, 8'd111}: color_data = 12'he00;
			{8'd114, 8'd112}: color_data = 12'he00;
			{8'd114, 8'd113}: color_data = 12'he00;
			{8'd114, 8'd114}: color_data = 12'he00;
			{8'd114, 8'd115}: color_data = 12'he00;
			{8'd114, 8'd116}: color_data = 12'he00;
			{8'd114, 8'd117}: color_data = 12'he00;
			{8'd114, 8'd118}: color_data = 12'he00;
			{8'd114, 8'd119}: color_data = 12'he00;
			{8'd114, 8'd120}: color_data = 12'he00;
			{8'd114, 8'd121}: color_data = 12'he00;
			{8'd114, 8'd122}: color_data = 12'he00;
			{8'd114, 8'd123}: color_data = 12'he00;
			{8'd114, 8'd124}: color_data = 12'he00;
			{8'd114, 8'd125}: color_data = 12'he00;
			{8'd114, 8'd126}: color_data = 12'he00;
			{8'd114, 8'd127}: color_data = 12'he00;
			{8'd114, 8'd128}: color_data = 12'he00;
			{8'd114, 8'd129}: color_data = 12'he00;
			{8'd114, 8'd130}: color_data = 12'he00;
			{8'd114, 8'd131}: color_data = 12'he00;
			{8'd114, 8'd132}: color_data = 12'he00;
			{8'd114, 8'd133}: color_data = 12'hf00;
			{8'd114, 8'd138}: color_data = 12'he00;
			{8'd114, 8'd139}: color_data = 12'he00;
			{8'd114, 8'd140}: color_data = 12'he00;
			{8'd114, 8'd141}: color_data = 12'he00;
			{8'd114, 8'd142}: color_data = 12'he00;
			{8'd114, 8'd143}: color_data = 12'he01;
			{8'd114, 8'd144}: color_data = 12'he00;
			{8'd115, 8'd4}: color_data = 12'h000;
			{8'd115, 8'd5}: color_data = 12'h000;
			{8'd115, 8'd6}: color_data = 12'h000;
			{8'd115, 8'd7}: color_data = 12'h392;
			{8'd115, 8'd8}: color_data = 12'h4b3;
			{8'd115, 8'd9}: color_data = 12'h4a3;
			{8'd115, 8'd10}: color_data = 12'h4a3;
			{8'd115, 8'd11}: color_data = 12'h4a3;
			{8'd115, 8'd12}: color_data = 12'h4b3;
			{8'd115, 8'd13}: color_data = 12'h261;
			{8'd115, 8'd14}: color_data = 12'h000;
			{8'd115, 8'd15}: color_data = 12'h000;
			{8'd115, 8'd16}: color_data = 12'h392;
			{8'd115, 8'd17}: color_data = 12'h392;
			{8'd115, 8'd18}: color_data = 12'h382;
			{8'd115, 8'd19}: color_data = 12'h272;
			{8'd115, 8'd20}: color_data = 12'h251;
			{8'd115, 8'd21}: color_data = 12'h010;
			{8'd115, 8'd22}: color_data = 12'h000;
			{8'd115, 8'd23}: color_data = 12'h130;
			{8'd115, 8'd24}: color_data = 12'h4b3;
			{8'd115, 8'd25}: color_data = 12'h4a3;
			{8'd115, 8'd26}: color_data = 12'h4a3;
			{8'd115, 8'd27}: color_data = 12'h4a3;
			{8'd115, 8'd28}: color_data = 12'h4a3;
			{8'd115, 8'd29}: color_data = 12'h4b3;
			{8'd115, 8'd30}: color_data = 12'h131;
			{8'd115, 8'd31}: color_data = 12'h000;
			{8'd115, 8'd32}: color_data = 12'h000;
			{8'd115, 8'd33}: color_data = 12'h000;
			{8'd115, 8'd34}: color_data = 12'h058;
			{8'd115, 8'd35}: color_data = 12'h0ae;
			{8'd115, 8'd36}: color_data = 12'h09d;
			{8'd115, 8'd37}: color_data = 12'h09d;
			{8'd115, 8'd38}: color_data = 12'h09d;
			{8'd115, 8'd39}: color_data = 12'h09d;
			{8'd115, 8'd40}: color_data = 12'h09d;
			{8'd115, 8'd41}: color_data = 12'h09d;
			{8'd115, 8'd42}: color_data = 12'h09d;
			{8'd115, 8'd43}: color_data = 12'h09d;
			{8'd115, 8'd44}: color_data = 12'h09d;
			{8'd115, 8'd45}: color_data = 12'h09d;
			{8'd115, 8'd46}: color_data = 12'h09d;
			{8'd115, 8'd47}: color_data = 12'h09d;
			{8'd115, 8'd48}: color_data = 12'h09d;
			{8'd115, 8'd49}: color_data = 12'h09d;
			{8'd115, 8'd50}: color_data = 12'h09d;
			{8'd115, 8'd51}: color_data = 12'h09d;
			{8'd115, 8'd52}: color_data = 12'h09d;
			{8'd115, 8'd53}: color_data = 12'h09d;
			{8'd115, 8'd54}: color_data = 12'h09d;
			{8'd115, 8'd55}: color_data = 12'h09d;
			{8'd115, 8'd56}: color_data = 12'h09d;
			{8'd115, 8'd57}: color_data = 12'h09d;
			{8'd115, 8'd58}: color_data = 12'h09d;
			{8'd115, 8'd59}: color_data = 12'h09d;
			{8'd115, 8'd60}: color_data = 12'h09d;
			{8'd115, 8'd61}: color_data = 12'h09d;
			{8'd115, 8'd62}: color_data = 12'h09d;
			{8'd115, 8'd63}: color_data = 12'h09d;
			{8'd115, 8'd64}: color_data = 12'h09d;
			{8'd115, 8'd65}: color_data = 12'h09d;
			{8'd115, 8'd66}: color_data = 12'h09d;
			{8'd115, 8'd67}: color_data = 12'h09c;
			{8'd115, 8'd68}: color_data = 12'h011;
			{8'd115, 8'd69}: color_data = 12'h000;
			{8'd115, 8'd70}: color_data = 12'h000;
			{8'd115, 8'd71}: color_data = 12'h000;
			{8'd115, 8'd72}: color_data = 12'h000;
			{8'd115, 8'd73}: color_data = 12'h000;
			{8'd115, 8'd74}: color_data = 12'h000;
			{8'd115, 8'd100}: color_data = 12'he00;
			{8'd115, 8'd101}: color_data = 12'hf01;
			{8'd115, 8'd102}: color_data = 12'he00;
			{8'd115, 8'd103}: color_data = 12'he00;
			{8'd115, 8'd104}: color_data = 12'he00;
			{8'd115, 8'd105}: color_data = 12'he00;
			{8'd115, 8'd106}: color_data = 12'hc00;
			{8'd115, 8'd111}: color_data = 12'he00;
			{8'd115, 8'd112}: color_data = 12'he01;
			{8'd115, 8'd113}: color_data = 12'hf01;
			{8'd115, 8'd114}: color_data = 12'he01;
			{8'd115, 8'd115}: color_data = 12'he01;
			{8'd115, 8'd116}: color_data = 12'he01;
			{8'd115, 8'd117}: color_data = 12'he01;
			{8'd115, 8'd118}: color_data = 12'he01;
			{8'd115, 8'd119}: color_data = 12'he00;
			{8'd115, 8'd120}: color_data = 12'he00;
			{8'd115, 8'd121}: color_data = 12'he00;
			{8'd115, 8'd122}: color_data = 12'he00;
			{8'd115, 8'd123}: color_data = 12'he00;
			{8'd115, 8'd124}: color_data = 12'he01;
			{8'd115, 8'd125}: color_data = 12'he00;
			{8'd115, 8'd126}: color_data = 12'he01;
			{8'd115, 8'd127}: color_data = 12'he01;
			{8'd115, 8'd128}: color_data = 12'he00;
			{8'd115, 8'd129}: color_data = 12'he00;
			{8'd115, 8'd130}: color_data = 12'he00;
			{8'd115, 8'd131}: color_data = 12'he00;
			{8'd115, 8'd132}: color_data = 12'he00;
			{8'd115, 8'd133}: color_data = 12'he00;
			{8'd115, 8'd138}: color_data = 12'he00;
			{8'd115, 8'd139}: color_data = 12'he00;
			{8'd115, 8'd140}: color_data = 12'he00;
			{8'd115, 8'd141}: color_data = 12'he00;
			{8'd115, 8'd142}: color_data = 12'he00;
			{8'd115, 8'd143}: color_data = 12'he01;
			{8'd115, 8'd144}: color_data = 12'he00;
			{8'd116, 8'd4}: color_data = 12'h000;
			{8'd116, 8'd5}: color_data = 12'h000;
			{8'd116, 8'd6}: color_data = 12'h000;
			{8'd116, 8'd7}: color_data = 12'h382;
			{8'd116, 8'd8}: color_data = 12'h4b3;
			{8'd116, 8'd9}: color_data = 12'h4a3;
			{8'd116, 8'd10}: color_data = 12'h4a3;
			{8'd116, 8'd11}: color_data = 12'h4a3;
			{8'd116, 8'd12}: color_data = 12'h4b3;
			{8'd116, 8'd13}: color_data = 12'h392;
			{8'd116, 8'd14}: color_data = 12'h000;
			{8'd116, 8'd15}: color_data = 12'h000;
			{8'd116, 8'd16}: color_data = 12'h000;
			{8'd116, 8'd17}: color_data = 12'h000;
			{8'd116, 8'd18}: color_data = 12'h000;
			{8'd116, 8'd19}: color_data = 12'h000;
			{8'd116, 8'd20}: color_data = 12'h000;
			{8'd116, 8'd21}: color_data = 12'h000;
			{8'd116, 8'd22}: color_data = 12'h000;
			{8'd116, 8'd23}: color_data = 12'h141;
			{8'd116, 8'd24}: color_data = 12'h4b3;
			{8'd116, 8'd25}: color_data = 12'h4b3;
			{8'd116, 8'd26}: color_data = 12'h4a3;
			{8'd116, 8'd27}: color_data = 12'h4a3;
			{8'd116, 8'd28}: color_data = 12'h4a3;
			{8'd116, 8'd29}: color_data = 12'h4b3;
			{8'd116, 8'd30}: color_data = 12'h131;
			{8'd116, 8'd31}: color_data = 12'h000;
			{8'd116, 8'd32}: color_data = 12'h000;
			{8'd116, 8'd33}: color_data = 12'h000;
			{8'd116, 8'd34}: color_data = 12'h034;
			{8'd116, 8'd35}: color_data = 12'h0ae;
			{8'd116, 8'd36}: color_data = 12'h09d;
			{8'd116, 8'd37}: color_data = 12'h09d;
			{8'd116, 8'd38}: color_data = 12'h09d;
			{8'd116, 8'd39}: color_data = 12'h09d;
			{8'd116, 8'd40}: color_data = 12'h09d;
			{8'd116, 8'd41}: color_data = 12'h09d;
			{8'd116, 8'd42}: color_data = 12'h09d;
			{8'd116, 8'd43}: color_data = 12'h09d;
			{8'd116, 8'd44}: color_data = 12'h09d;
			{8'd116, 8'd45}: color_data = 12'h09d;
			{8'd116, 8'd46}: color_data = 12'h09d;
			{8'd116, 8'd47}: color_data = 12'h09d;
			{8'd116, 8'd48}: color_data = 12'h09d;
			{8'd116, 8'd49}: color_data = 12'h09d;
			{8'd116, 8'd50}: color_data = 12'h09d;
			{8'd116, 8'd51}: color_data = 12'h09d;
			{8'd116, 8'd52}: color_data = 12'h09d;
			{8'd116, 8'd53}: color_data = 12'h09d;
			{8'd116, 8'd54}: color_data = 12'h09d;
			{8'd116, 8'd55}: color_data = 12'h09d;
			{8'd116, 8'd56}: color_data = 12'h09d;
			{8'd116, 8'd57}: color_data = 12'h09d;
			{8'd116, 8'd58}: color_data = 12'h09d;
			{8'd116, 8'd59}: color_data = 12'h09d;
			{8'd116, 8'd60}: color_data = 12'h09d;
			{8'd116, 8'd61}: color_data = 12'h09d;
			{8'd116, 8'd62}: color_data = 12'h09d;
			{8'd116, 8'd63}: color_data = 12'h09d;
			{8'd116, 8'd64}: color_data = 12'h09d;
			{8'd116, 8'd65}: color_data = 12'h09d;
			{8'd116, 8'd66}: color_data = 12'h09d;
			{8'd116, 8'd67}: color_data = 12'h08c;
			{8'd116, 8'd68}: color_data = 12'h001;
			{8'd116, 8'd69}: color_data = 12'h000;
			{8'd116, 8'd70}: color_data = 12'h000;
			{8'd116, 8'd71}: color_data = 12'h000;
			{8'd116, 8'd72}: color_data = 12'h000;
			{8'd116, 8'd73}: color_data = 12'h000;
			{8'd116, 8'd74}: color_data = 12'h000;
			{8'd116, 8'd100}: color_data = 12'he00;
			{8'd116, 8'd101}: color_data = 12'hf01;
			{8'd116, 8'd102}: color_data = 12'he00;
			{8'd116, 8'd103}: color_data = 12'he00;
			{8'd116, 8'd104}: color_data = 12'he00;
			{8'd116, 8'd105}: color_data = 12'he00;
			{8'd116, 8'd106}: color_data = 12'hc00;
			{8'd116, 8'd111}: color_data = 12'he01;
			{8'd116, 8'd112}: color_data = 12'he00;
			{8'd116, 8'd113}: color_data = 12'he00;
			{8'd116, 8'd114}: color_data = 12'he00;
			{8'd116, 8'd115}: color_data = 12'he00;
			{8'd116, 8'd116}: color_data = 12'he00;
			{8'd116, 8'd117}: color_data = 12'he00;
			{8'd116, 8'd118}: color_data = 12'he00;
			{8'd116, 8'd119}: color_data = 12'he00;
			{8'd116, 8'd120}: color_data = 12'he00;
			{8'd116, 8'd121}: color_data = 12'he00;
			{8'd116, 8'd122}: color_data = 12'he00;
			{8'd116, 8'd123}: color_data = 12'he00;
			{8'd116, 8'd124}: color_data = 12'he00;
			{8'd116, 8'd125}: color_data = 12'he00;
			{8'd116, 8'd126}: color_data = 12'he00;
			{8'd116, 8'd127}: color_data = 12'he00;
			{8'd116, 8'd128}: color_data = 12'he00;
			{8'd116, 8'd129}: color_data = 12'he00;
			{8'd116, 8'd130}: color_data = 12'he00;
			{8'd116, 8'd131}: color_data = 12'he00;
			{8'd116, 8'd132}: color_data = 12'hf01;
			{8'd116, 8'd133}: color_data = 12'he00;
			{8'd116, 8'd138}: color_data = 12'he00;
			{8'd116, 8'd139}: color_data = 12'he00;
			{8'd116, 8'd140}: color_data = 12'he00;
			{8'd116, 8'd141}: color_data = 12'he00;
			{8'd116, 8'd142}: color_data = 12'he00;
			{8'd116, 8'd143}: color_data = 12'he01;
			{8'd116, 8'd144}: color_data = 12'he00;
			{8'd117, 8'd3}: color_data = 12'h000;
			{8'd117, 8'd4}: color_data = 12'h000;
			{8'd117, 8'd5}: color_data = 12'h000;
			{8'd117, 8'd6}: color_data = 12'h000;
			{8'd117, 8'd7}: color_data = 12'h261;
			{8'd117, 8'd8}: color_data = 12'h4b3;
			{8'd117, 8'd9}: color_data = 12'h4b3;
			{8'd117, 8'd10}: color_data = 12'h4b3;
			{8'd117, 8'd11}: color_data = 12'h4b3;
			{8'd117, 8'd12}: color_data = 12'h4b3;
			{8'd117, 8'd13}: color_data = 12'h4a3;
			{8'd117, 8'd14}: color_data = 12'h010;
			{8'd117, 8'd15}: color_data = 12'h000;
			{8'd117, 8'd16}: color_data = 12'h000;
			{8'd117, 8'd17}: color_data = 12'h000;
			{8'd117, 8'd18}: color_data = 12'h000;
			{8'd117, 8'd19}: color_data = 12'h000;
			{8'd117, 8'd20}: color_data = 12'h000;
			{8'd117, 8'd21}: color_data = 12'h000;
			{8'd117, 8'd22}: color_data = 12'h000;
			{8'd117, 8'd23}: color_data = 12'h141;
			{8'd117, 8'd24}: color_data = 12'h3a3;
			{8'd117, 8'd25}: color_data = 12'h4a3;
			{8'd117, 8'd26}: color_data = 12'h4b3;
			{8'd117, 8'd27}: color_data = 12'h4b3;
			{8'd117, 8'd28}: color_data = 12'h4b3;
			{8'd117, 8'd29}: color_data = 12'h4b3;
			{8'd117, 8'd30}: color_data = 12'h141;
			{8'd117, 8'd31}: color_data = 12'h000;
			{8'd117, 8'd32}: color_data = 12'h000;
			{8'd117, 8'd33}: color_data = 12'h000;
			{8'd117, 8'd34}: color_data = 12'h012;
			{8'd117, 8'd35}: color_data = 12'h09d;
			{8'd117, 8'd36}: color_data = 12'h09d;
			{8'd117, 8'd37}: color_data = 12'h09d;
			{8'd117, 8'd38}: color_data = 12'h09d;
			{8'd117, 8'd39}: color_data = 12'h09d;
			{8'd117, 8'd40}: color_data = 12'h09d;
			{8'd117, 8'd41}: color_data = 12'h09d;
			{8'd117, 8'd42}: color_data = 12'h09d;
			{8'd117, 8'd43}: color_data = 12'h09d;
			{8'd117, 8'd44}: color_data = 12'h09d;
			{8'd117, 8'd45}: color_data = 12'h09d;
			{8'd117, 8'd46}: color_data = 12'h09d;
			{8'd117, 8'd47}: color_data = 12'h09d;
			{8'd117, 8'd48}: color_data = 12'h09d;
			{8'd117, 8'd49}: color_data = 12'h09d;
			{8'd117, 8'd50}: color_data = 12'h09d;
			{8'd117, 8'd51}: color_data = 12'h09d;
			{8'd117, 8'd52}: color_data = 12'h09d;
			{8'd117, 8'd53}: color_data = 12'h09d;
			{8'd117, 8'd54}: color_data = 12'h09d;
			{8'd117, 8'd55}: color_data = 12'h09d;
			{8'd117, 8'd56}: color_data = 12'h09d;
			{8'd117, 8'd57}: color_data = 12'h09d;
			{8'd117, 8'd58}: color_data = 12'h09d;
			{8'd117, 8'd59}: color_data = 12'h09d;
			{8'd117, 8'd60}: color_data = 12'h09d;
			{8'd117, 8'd61}: color_data = 12'h09d;
			{8'd117, 8'd62}: color_data = 12'h09d;
			{8'd117, 8'd63}: color_data = 12'h09d;
			{8'd117, 8'd64}: color_data = 12'h09d;
			{8'd117, 8'd65}: color_data = 12'h09d;
			{8'd117, 8'd66}: color_data = 12'h09d;
			{8'd117, 8'd67}: color_data = 12'h08b;
			{8'd117, 8'd68}: color_data = 12'h000;
			{8'd117, 8'd69}: color_data = 12'h000;
			{8'd117, 8'd70}: color_data = 12'h000;
			{8'd117, 8'd71}: color_data = 12'h000;
			{8'd117, 8'd72}: color_data = 12'h000;
			{8'd117, 8'd73}: color_data = 12'h000;
			{8'd117, 8'd74}: color_data = 12'h000;
			{8'd117, 8'd100}: color_data = 12'he00;
			{8'd117, 8'd101}: color_data = 12'hf01;
			{8'd117, 8'd102}: color_data = 12'he00;
			{8'd117, 8'd103}: color_data = 12'he00;
			{8'd117, 8'd104}: color_data = 12'he00;
			{8'd117, 8'd105}: color_data = 12'he00;
			{8'd117, 8'd106}: color_data = 12'hc00;
			{8'd117, 8'd111}: color_data = 12'he01;
			{8'd117, 8'd112}: color_data = 12'he00;
			{8'd117, 8'd113}: color_data = 12'he00;
			{8'd117, 8'd114}: color_data = 12'he00;
			{8'd117, 8'd115}: color_data = 12'he00;
			{8'd117, 8'd116}: color_data = 12'he00;
			{8'd117, 8'd117}: color_data = 12'he00;
			{8'd117, 8'd118}: color_data = 12'he00;
			{8'd117, 8'd119}: color_data = 12'he00;
			{8'd117, 8'd120}: color_data = 12'he00;
			{8'd117, 8'd121}: color_data = 12'he00;
			{8'd117, 8'd122}: color_data = 12'he00;
			{8'd117, 8'd123}: color_data = 12'he00;
			{8'd117, 8'd124}: color_data = 12'he00;
			{8'd117, 8'd125}: color_data = 12'he00;
			{8'd117, 8'd126}: color_data = 12'he00;
			{8'd117, 8'd127}: color_data = 12'he00;
			{8'd117, 8'd128}: color_data = 12'he00;
			{8'd117, 8'd129}: color_data = 12'he00;
			{8'd117, 8'd130}: color_data = 12'he00;
			{8'd117, 8'd131}: color_data = 12'he00;
			{8'd117, 8'd132}: color_data = 12'hf01;
			{8'd117, 8'd133}: color_data = 12'he00;
			{8'd117, 8'd138}: color_data = 12'he00;
			{8'd117, 8'd139}: color_data = 12'he00;
			{8'd117, 8'd140}: color_data = 12'he00;
			{8'd117, 8'd141}: color_data = 12'he00;
			{8'd117, 8'd142}: color_data = 12'he00;
			{8'd117, 8'd143}: color_data = 12'he01;
			{8'd117, 8'd144}: color_data = 12'he00;
			{8'd118, 8'd3}: color_data = 12'h000;
			{8'd118, 8'd4}: color_data = 12'h000;
			{8'd118, 8'd5}: color_data = 12'h000;
			{8'd118, 8'd6}: color_data = 12'h000;
			{8'd118, 8'd7}: color_data = 12'h141;
			{8'd118, 8'd8}: color_data = 12'h4a3;
			{8'd118, 8'd9}: color_data = 12'h392;
			{8'd118, 8'd10}: color_data = 12'h372;
			{8'd118, 8'd11}: color_data = 12'h251;
			{8'd118, 8'd12}: color_data = 12'h141;
			{8'd118, 8'd13}: color_data = 12'h120;
			{8'd118, 8'd14}: color_data = 12'h000;
			{8'd118, 8'd15}: color_data = 12'h000;
			{8'd118, 8'd16}: color_data = 12'h000;
			{8'd118, 8'd17}: color_data = 12'h000;
			{8'd118, 8'd18}: color_data = 12'h000;
			{8'd118, 8'd19}: color_data = 12'h000;
			{8'd118, 8'd20}: color_data = 12'h000;
			{8'd118, 8'd21}: color_data = 12'h000;
			{8'd118, 8'd22}: color_data = 12'h000;
			{8'd118, 8'd23}: color_data = 12'h000;
			{8'd118, 8'd24}: color_data = 12'h000;
			{8'd118, 8'd25}: color_data = 12'h010;
			{8'd118, 8'd26}: color_data = 12'h130;
			{8'd118, 8'd27}: color_data = 12'h141;
			{8'd118, 8'd28}: color_data = 12'h261;
			{8'd118, 8'd29}: color_data = 12'h382;
			{8'd118, 8'd30}: color_data = 12'h131;
			{8'd118, 8'd31}: color_data = 12'h000;
			{8'd118, 8'd32}: color_data = 12'h000;
			{8'd118, 8'd33}: color_data = 12'h000;
			{8'd118, 8'd34}: color_data = 12'h000;
			{8'd118, 8'd35}: color_data = 12'h08b;
			{8'd118, 8'd36}: color_data = 12'h09d;
			{8'd118, 8'd37}: color_data = 12'h09d;
			{8'd118, 8'd38}: color_data = 12'h09d;
			{8'd118, 8'd39}: color_data = 12'h09d;
			{8'd118, 8'd40}: color_data = 12'h09d;
			{8'd118, 8'd41}: color_data = 12'h09d;
			{8'd118, 8'd42}: color_data = 12'h09d;
			{8'd118, 8'd43}: color_data = 12'h09d;
			{8'd118, 8'd44}: color_data = 12'h09d;
			{8'd118, 8'd45}: color_data = 12'h09d;
			{8'd118, 8'd46}: color_data = 12'h09d;
			{8'd118, 8'd47}: color_data = 12'h09d;
			{8'd118, 8'd48}: color_data = 12'h09d;
			{8'd118, 8'd49}: color_data = 12'h09d;
			{8'd118, 8'd50}: color_data = 12'h09d;
			{8'd118, 8'd51}: color_data = 12'h09d;
			{8'd118, 8'd52}: color_data = 12'h09d;
			{8'd118, 8'd53}: color_data = 12'h09d;
			{8'd118, 8'd54}: color_data = 12'h09d;
			{8'd118, 8'd55}: color_data = 12'h09d;
			{8'd118, 8'd56}: color_data = 12'h09d;
			{8'd118, 8'd57}: color_data = 12'h09d;
			{8'd118, 8'd58}: color_data = 12'h09d;
			{8'd118, 8'd59}: color_data = 12'h09d;
			{8'd118, 8'd60}: color_data = 12'h09d;
			{8'd118, 8'd61}: color_data = 12'h09d;
			{8'd118, 8'd62}: color_data = 12'h09d;
			{8'd118, 8'd63}: color_data = 12'h09d;
			{8'd118, 8'd64}: color_data = 12'h09d;
			{8'd118, 8'd65}: color_data = 12'h09d;
			{8'd118, 8'd66}: color_data = 12'h09d;
			{8'd118, 8'd67}: color_data = 12'h07b;
			{8'd118, 8'd68}: color_data = 12'h000;
			{8'd118, 8'd69}: color_data = 12'h000;
			{8'd118, 8'd70}: color_data = 12'h000;
			{8'd118, 8'd71}: color_data = 12'h000;
			{8'd118, 8'd72}: color_data = 12'h000;
			{8'd118, 8'd73}: color_data = 12'h000;
			{8'd118, 8'd74}: color_data = 12'h000;
			{8'd118, 8'd100}: color_data = 12'he00;
			{8'd118, 8'd101}: color_data = 12'hf01;
			{8'd118, 8'd102}: color_data = 12'he00;
			{8'd118, 8'd103}: color_data = 12'he00;
			{8'd118, 8'd104}: color_data = 12'he00;
			{8'd118, 8'd105}: color_data = 12'he00;
			{8'd118, 8'd106}: color_data = 12'hc00;
			{8'd118, 8'd111}: color_data = 12'he01;
			{8'd118, 8'd112}: color_data = 12'he00;
			{8'd118, 8'd113}: color_data = 12'he00;
			{8'd118, 8'd114}: color_data = 12'he00;
			{8'd118, 8'd115}: color_data = 12'he00;
			{8'd118, 8'd116}: color_data = 12'he00;
			{8'd118, 8'd117}: color_data = 12'he00;
			{8'd118, 8'd118}: color_data = 12'he00;
			{8'd118, 8'd119}: color_data = 12'he00;
			{8'd118, 8'd120}: color_data = 12'he00;
			{8'd118, 8'd121}: color_data = 12'he00;
			{8'd118, 8'd122}: color_data = 12'he00;
			{8'd118, 8'd123}: color_data = 12'he00;
			{8'd118, 8'd124}: color_data = 12'he00;
			{8'd118, 8'd125}: color_data = 12'he00;
			{8'd118, 8'd126}: color_data = 12'he00;
			{8'd118, 8'd127}: color_data = 12'he00;
			{8'd118, 8'd128}: color_data = 12'he00;
			{8'd118, 8'd129}: color_data = 12'he00;
			{8'd118, 8'd130}: color_data = 12'he00;
			{8'd118, 8'd131}: color_data = 12'he00;
			{8'd118, 8'd132}: color_data = 12'hf01;
			{8'd118, 8'd133}: color_data = 12'he00;
			{8'd118, 8'd138}: color_data = 12'he00;
			{8'd118, 8'd139}: color_data = 12'he00;
			{8'd118, 8'd140}: color_data = 12'he00;
			{8'd118, 8'd141}: color_data = 12'he00;
			{8'd118, 8'd142}: color_data = 12'he00;
			{8'd118, 8'd143}: color_data = 12'he01;
			{8'd118, 8'd144}: color_data = 12'he00;
			{8'd119, 8'd3}: color_data = 12'h000;
			{8'd119, 8'd4}: color_data = 12'h000;
			{8'd119, 8'd5}: color_data = 12'h000;
			{8'd119, 8'd6}: color_data = 12'h000;
			{8'd119, 8'd7}: color_data = 12'h000;
			{8'd119, 8'd8}: color_data = 12'h010;
			{8'd119, 8'd9}: color_data = 12'h000;
			{8'd119, 8'd10}: color_data = 12'h000;
			{8'd119, 8'd11}: color_data = 12'h000;
			{8'd119, 8'd12}: color_data = 12'h000;
			{8'd119, 8'd13}: color_data = 12'h000;
			{8'd119, 8'd14}: color_data = 12'h000;
			{8'd119, 8'd15}: color_data = 12'h000;
			{8'd119, 8'd16}: color_data = 12'h000;
			{8'd119, 8'd17}: color_data = 12'h000;
			{8'd119, 8'd18}: color_data = 12'h000;
			{8'd119, 8'd19}: color_data = 12'h000;
			{8'd119, 8'd20}: color_data = 12'h000;
			{8'd119, 8'd21}: color_data = 12'h000;
			{8'd119, 8'd22}: color_data = 12'h000;
			{8'd119, 8'd23}: color_data = 12'h000;
			{8'd119, 8'd24}: color_data = 12'h000;
			{8'd119, 8'd25}: color_data = 12'h000;
			{8'd119, 8'd26}: color_data = 12'h000;
			{8'd119, 8'd27}: color_data = 12'h000;
			{8'd119, 8'd28}: color_data = 12'h000;
			{8'd119, 8'd29}: color_data = 12'h000;
			{8'd119, 8'd30}: color_data = 12'h000;
			{8'd119, 8'd31}: color_data = 12'h000;
			{8'd119, 8'd32}: color_data = 12'h000;
			{8'd119, 8'd33}: color_data = 12'h000;
			{8'd119, 8'd34}: color_data = 12'h000;
			{8'd119, 8'd35}: color_data = 12'h068;
			{8'd119, 8'd36}: color_data = 12'h0ae;
			{8'd119, 8'd37}: color_data = 12'h09d;
			{8'd119, 8'd38}: color_data = 12'h09d;
			{8'd119, 8'd39}: color_data = 12'h09d;
			{8'd119, 8'd40}: color_data = 12'h09d;
			{8'd119, 8'd41}: color_data = 12'h09d;
			{8'd119, 8'd42}: color_data = 12'h09d;
			{8'd119, 8'd43}: color_data = 12'h09d;
			{8'd119, 8'd44}: color_data = 12'h09d;
			{8'd119, 8'd45}: color_data = 12'h09d;
			{8'd119, 8'd46}: color_data = 12'h09d;
			{8'd119, 8'd47}: color_data = 12'h09d;
			{8'd119, 8'd48}: color_data = 12'h09d;
			{8'd119, 8'd49}: color_data = 12'h09d;
			{8'd119, 8'd50}: color_data = 12'h09d;
			{8'd119, 8'd51}: color_data = 12'h09d;
			{8'd119, 8'd52}: color_data = 12'h09d;
			{8'd119, 8'd53}: color_data = 12'h09d;
			{8'd119, 8'd54}: color_data = 12'h09d;
			{8'd119, 8'd55}: color_data = 12'h09d;
			{8'd119, 8'd56}: color_data = 12'h09d;
			{8'd119, 8'd57}: color_data = 12'h09d;
			{8'd119, 8'd58}: color_data = 12'h09d;
			{8'd119, 8'd59}: color_data = 12'h09d;
			{8'd119, 8'd60}: color_data = 12'h09d;
			{8'd119, 8'd61}: color_data = 12'h09d;
			{8'd119, 8'd62}: color_data = 12'h09d;
			{8'd119, 8'd63}: color_data = 12'h09d;
			{8'd119, 8'd64}: color_data = 12'h09d;
			{8'd119, 8'd65}: color_data = 12'h09d;
			{8'd119, 8'd66}: color_data = 12'h0ae;
			{8'd119, 8'd67}: color_data = 12'h07a;
			{8'd119, 8'd68}: color_data = 12'h000;
			{8'd119, 8'd69}: color_data = 12'h000;
			{8'd119, 8'd70}: color_data = 12'h000;
			{8'd119, 8'd71}: color_data = 12'h000;
			{8'd119, 8'd72}: color_data = 12'h000;
			{8'd119, 8'd73}: color_data = 12'h000;
			{8'd119, 8'd74}: color_data = 12'h000;
			{8'd119, 8'd100}: color_data = 12'he00;
			{8'd119, 8'd101}: color_data = 12'hf01;
			{8'd119, 8'd102}: color_data = 12'he00;
			{8'd119, 8'd103}: color_data = 12'he00;
			{8'd119, 8'd104}: color_data = 12'he00;
			{8'd119, 8'd105}: color_data = 12'he00;
			{8'd119, 8'd106}: color_data = 12'hc00;
			{8'd119, 8'd111}: color_data = 12'he00;
			{8'd119, 8'd112}: color_data = 12'he00;
			{8'd119, 8'd113}: color_data = 12'he00;
			{8'd119, 8'd114}: color_data = 12'he00;
			{8'd119, 8'd115}: color_data = 12'he00;
			{8'd119, 8'd116}: color_data = 12'he00;
			{8'd119, 8'd117}: color_data = 12'he00;
			{8'd119, 8'd118}: color_data = 12'he00;
			{8'd119, 8'd119}: color_data = 12'he00;
			{8'd119, 8'd120}: color_data = 12'he00;
			{8'd119, 8'd121}: color_data = 12'he00;
			{8'd119, 8'd122}: color_data = 12'he00;
			{8'd119, 8'd123}: color_data = 12'he00;
			{8'd119, 8'd124}: color_data = 12'he00;
			{8'd119, 8'd125}: color_data = 12'he00;
			{8'd119, 8'd126}: color_data = 12'he00;
			{8'd119, 8'd127}: color_data = 12'he00;
			{8'd119, 8'd128}: color_data = 12'he00;
			{8'd119, 8'd129}: color_data = 12'he00;
			{8'd119, 8'd130}: color_data = 12'he00;
			{8'd119, 8'd131}: color_data = 12'he00;
			{8'd119, 8'd132}: color_data = 12'hf01;
			{8'd119, 8'd133}: color_data = 12'he00;
			{8'd119, 8'd138}: color_data = 12'he00;
			{8'd119, 8'd139}: color_data = 12'he00;
			{8'd119, 8'd140}: color_data = 12'he00;
			{8'd119, 8'd141}: color_data = 12'he00;
			{8'd119, 8'd142}: color_data = 12'he00;
			{8'd119, 8'd143}: color_data = 12'he01;
			{8'd119, 8'd144}: color_data = 12'he00;
			{8'd120, 8'd2}: color_data = 12'h000;
			{8'd120, 8'd3}: color_data = 12'h000;
			{8'd120, 8'd4}: color_data = 12'h000;
			{8'd120, 8'd5}: color_data = 12'h440;
			{8'd120, 8'd6}: color_data = 12'h000;
			{8'd120, 8'd7}: color_data = 12'h000;
			{8'd120, 8'd8}: color_data = 12'h000;
			{8'd120, 8'd9}: color_data = 12'h000;
			{8'd120, 8'd10}: color_data = 12'h110;
			{8'd120, 8'd11}: color_data = 12'h320;
			{8'd120, 8'd12}: color_data = 12'h540;
			{8'd120, 8'd13}: color_data = 12'h860;
			{8'd120, 8'd14}: color_data = 12'h970;
			{8'd120, 8'd15}: color_data = 12'h760;
			{8'd120, 8'd16}: color_data = 12'h540;
			{8'd120, 8'd17}: color_data = 12'h430;
			{8'd120, 8'd18}: color_data = 12'h320;
			{8'd120, 8'd19}: color_data = 12'h110;
			{8'd120, 8'd20}: color_data = 12'h000;
			{8'd120, 8'd21}: color_data = 12'h000;
			{8'd120, 8'd22}: color_data = 12'h000;
			{8'd120, 8'd23}: color_data = 12'h000;
			{8'd120, 8'd24}: color_data = 12'h000;
			{8'd120, 8'd25}: color_data = 12'h000;
			{8'd120, 8'd26}: color_data = 12'h000;
			{8'd120, 8'd27}: color_data = 12'h000;
			{8'd120, 8'd28}: color_data = 12'h000;
			{8'd120, 8'd29}: color_data = 12'h000;
			{8'd120, 8'd30}: color_data = 12'h000;
			{8'd120, 8'd31}: color_data = 12'h000;
			{8'd120, 8'd32}: color_data = 12'h000;
			{8'd120, 8'd33}: color_data = 12'h000;
			{8'd120, 8'd34}: color_data = 12'h000;
			{8'd120, 8'd35}: color_data = 12'h035;
			{8'd120, 8'd36}: color_data = 12'h0ae;
			{8'd120, 8'd37}: color_data = 12'h09d;
			{8'd120, 8'd38}: color_data = 12'h09d;
			{8'd120, 8'd39}: color_data = 12'h09d;
			{8'd120, 8'd40}: color_data = 12'h09d;
			{8'd120, 8'd41}: color_data = 12'h09d;
			{8'd120, 8'd42}: color_data = 12'h09d;
			{8'd120, 8'd43}: color_data = 12'h09d;
			{8'd120, 8'd44}: color_data = 12'h09d;
			{8'd120, 8'd45}: color_data = 12'h09d;
			{8'd120, 8'd46}: color_data = 12'h09d;
			{8'd120, 8'd47}: color_data = 12'h09d;
			{8'd120, 8'd48}: color_data = 12'h09d;
			{8'd120, 8'd49}: color_data = 12'h09d;
			{8'd120, 8'd50}: color_data = 12'h09d;
			{8'd120, 8'd51}: color_data = 12'h09d;
			{8'd120, 8'd52}: color_data = 12'h09d;
			{8'd120, 8'd53}: color_data = 12'h09d;
			{8'd120, 8'd54}: color_data = 12'h09d;
			{8'd120, 8'd55}: color_data = 12'h09d;
			{8'd120, 8'd56}: color_data = 12'h09d;
			{8'd120, 8'd57}: color_data = 12'h09d;
			{8'd120, 8'd58}: color_data = 12'h09d;
			{8'd120, 8'd59}: color_data = 12'h09d;
			{8'd120, 8'd60}: color_data = 12'h09d;
			{8'd120, 8'd61}: color_data = 12'h0ae;
			{8'd120, 8'd62}: color_data = 12'h0ae;
			{8'd120, 8'd63}: color_data = 12'h0ae;
			{8'd120, 8'd64}: color_data = 12'h09d;
			{8'd120, 8'd65}: color_data = 12'h08c;
			{8'd120, 8'd66}: color_data = 12'h07a;
			{8'd120, 8'd67}: color_data = 12'h045;
			{8'd120, 8'd68}: color_data = 12'h000;
			{8'd120, 8'd69}: color_data = 12'h000;
			{8'd120, 8'd70}: color_data = 12'h000;
			{8'd120, 8'd71}: color_data = 12'h000;
			{8'd120, 8'd72}: color_data = 12'h000;
			{8'd120, 8'd73}: color_data = 12'h000;
			{8'd120, 8'd74}: color_data = 12'h000;
			{8'd120, 8'd100}: color_data = 12'he00;
			{8'd120, 8'd101}: color_data = 12'hf01;
			{8'd120, 8'd102}: color_data = 12'he00;
			{8'd120, 8'd103}: color_data = 12'he00;
			{8'd120, 8'd104}: color_data = 12'he00;
			{8'd120, 8'd105}: color_data = 12'he00;
			{8'd120, 8'd106}: color_data = 12'hc00;
			{8'd120, 8'd111}: color_data = 12'he00;
			{8'd120, 8'd112}: color_data = 12'he00;
			{8'd120, 8'd113}: color_data = 12'he00;
			{8'd120, 8'd114}: color_data = 12'he00;
			{8'd120, 8'd115}: color_data = 12'he00;
			{8'd120, 8'd116}: color_data = 12'he00;
			{8'd120, 8'd117}: color_data = 12'he00;
			{8'd120, 8'd118}: color_data = 12'he00;
			{8'd120, 8'd119}: color_data = 12'he00;
			{8'd120, 8'd120}: color_data = 12'he00;
			{8'd120, 8'd121}: color_data = 12'he00;
			{8'd120, 8'd122}: color_data = 12'he00;
			{8'd120, 8'd123}: color_data = 12'he00;
			{8'd120, 8'd124}: color_data = 12'he00;
			{8'd120, 8'd125}: color_data = 12'he00;
			{8'd120, 8'd126}: color_data = 12'he00;
			{8'd120, 8'd127}: color_data = 12'he00;
			{8'd120, 8'd128}: color_data = 12'he00;
			{8'd120, 8'd129}: color_data = 12'he00;
			{8'd120, 8'd130}: color_data = 12'he00;
			{8'd120, 8'd131}: color_data = 12'he00;
			{8'd120, 8'd132}: color_data = 12'he00;
			{8'd120, 8'd133}: color_data = 12'he00;
			{8'd120, 8'd138}: color_data = 12'he00;
			{8'd120, 8'd139}: color_data = 12'he00;
			{8'd120, 8'd140}: color_data = 12'he00;
			{8'd120, 8'd141}: color_data = 12'he00;
			{8'd120, 8'd142}: color_data = 12'he00;
			{8'd120, 8'd143}: color_data = 12'he01;
			{8'd120, 8'd144}: color_data = 12'he00;
			{8'd121, 8'd2}: color_data = 12'h000;
			{8'd121, 8'd3}: color_data = 12'h000;
			{8'd121, 8'd4}: color_data = 12'h000;
			{8'd121, 8'd5}: color_data = 12'ha80;
			{8'd121, 8'd6}: color_data = 12'h650;
			{8'd121, 8'd7}: color_data = 12'h760;
			{8'd121, 8'd8}: color_data = 12'ha80;
			{8'd121, 8'd9}: color_data = 12'hca0;
			{8'd121, 8'd10}: color_data = 12'hec0;
			{8'd121, 8'd11}: color_data = 12'hfc0;
			{8'd121, 8'd12}: color_data = 12'hfd0;
			{8'd121, 8'd13}: color_data = 12'hfd0;
			{8'd121, 8'd14}: color_data = 12'hfd0;
			{8'd121, 8'd15}: color_data = 12'hfd0;
			{8'd121, 8'd16}: color_data = 12'hfd0;
			{8'd121, 8'd17}: color_data = 12'hfd0;
			{8'd121, 8'd18}: color_data = 12'hfc0;
			{8'd121, 8'd19}: color_data = 12'hec0;
			{8'd121, 8'd20}: color_data = 12'hdb0;
			{8'd121, 8'd21}: color_data = 12'hca0;
			{8'd121, 8'd22}: color_data = 12'hb90;
			{8'd121, 8'd23}: color_data = 12'ha80;
			{8'd121, 8'd24}: color_data = 12'h870;
			{8'd121, 8'd25}: color_data = 12'h650;
			{8'd121, 8'd26}: color_data = 12'h540;
			{8'd121, 8'd27}: color_data = 12'h430;
			{8'd121, 8'd28}: color_data = 12'h220;
			{8'd121, 8'd29}: color_data = 12'h110;
			{8'd121, 8'd30}: color_data = 12'h000;
			{8'd121, 8'd31}: color_data = 12'h000;
			{8'd121, 8'd32}: color_data = 12'h000;
			{8'd121, 8'd33}: color_data = 12'h000;
			{8'd121, 8'd34}: color_data = 12'h000;
			{8'd121, 8'd35}: color_data = 12'h012;
			{8'd121, 8'd36}: color_data = 12'h09d;
			{8'd121, 8'd37}: color_data = 12'h09d;
			{8'd121, 8'd38}: color_data = 12'h09d;
			{8'd121, 8'd39}: color_data = 12'h09d;
			{8'd121, 8'd40}: color_data = 12'h09d;
			{8'd121, 8'd41}: color_data = 12'h09d;
			{8'd121, 8'd42}: color_data = 12'h09d;
			{8'd121, 8'd43}: color_data = 12'h09d;
			{8'd121, 8'd44}: color_data = 12'h09d;
			{8'd121, 8'd45}: color_data = 12'h09d;
			{8'd121, 8'd46}: color_data = 12'h09d;
			{8'd121, 8'd47}: color_data = 12'h09d;
			{8'd121, 8'd48}: color_data = 12'h09d;
			{8'd121, 8'd49}: color_data = 12'h09d;
			{8'd121, 8'd50}: color_data = 12'h09d;
			{8'd121, 8'd51}: color_data = 12'h09d;
			{8'd121, 8'd52}: color_data = 12'h09d;
			{8'd121, 8'd53}: color_data = 12'h09d;
			{8'd121, 8'd54}: color_data = 12'h09d;
			{8'd121, 8'd55}: color_data = 12'h09d;
			{8'd121, 8'd56}: color_data = 12'h0ae;
			{8'd121, 8'd57}: color_data = 12'h0ae;
			{8'd121, 8'd58}: color_data = 12'h09d;
			{8'd121, 8'd59}: color_data = 12'h09c;
			{8'd121, 8'd60}: color_data = 12'h08b;
			{8'd121, 8'd61}: color_data = 12'h069;
			{8'd121, 8'd62}: color_data = 12'h057;
			{8'd121, 8'd63}: color_data = 12'h034;
			{8'd121, 8'd64}: color_data = 12'h012;
			{8'd121, 8'd65}: color_data = 12'h001;
			{8'd121, 8'd66}: color_data = 12'h000;
			{8'd121, 8'd67}: color_data = 12'h000;
			{8'd121, 8'd68}: color_data = 12'h000;
			{8'd121, 8'd69}: color_data = 12'h000;
			{8'd121, 8'd70}: color_data = 12'h000;
			{8'd121, 8'd71}: color_data = 12'h000;
			{8'd121, 8'd72}: color_data = 12'h000;
			{8'd121, 8'd73}: color_data = 12'h000;
			{8'd121, 8'd74}: color_data = 12'h000;
			{8'd121, 8'd100}: color_data = 12'he00;
			{8'd121, 8'd101}: color_data = 12'hf01;
			{8'd121, 8'd102}: color_data = 12'he00;
			{8'd121, 8'd103}: color_data = 12'he00;
			{8'd121, 8'd104}: color_data = 12'he00;
			{8'd121, 8'd105}: color_data = 12'he00;
			{8'd121, 8'd106}: color_data = 12'hc00;
			{8'd121, 8'd138}: color_data = 12'he00;
			{8'd121, 8'd139}: color_data = 12'he00;
			{8'd121, 8'd140}: color_data = 12'he00;
			{8'd121, 8'd141}: color_data = 12'he00;
			{8'd121, 8'd142}: color_data = 12'he00;
			{8'd121, 8'd143}: color_data = 12'he01;
			{8'd121, 8'd144}: color_data = 12'he00;
			{8'd122, 8'd2}: color_data = 12'h000;
			{8'd122, 8'd3}: color_data = 12'h000;
			{8'd122, 8'd4}: color_data = 12'h100;
			{8'd122, 8'd5}: color_data = 12'heb0;
			{8'd122, 8'd6}: color_data = 12'hfd0;
			{8'd122, 8'd7}: color_data = 12'hfd0;
			{8'd122, 8'd8}: color_data = 12'hfd0;
			{8'd122, 8'd9}: color_data = 12'hfd0;
			{8'd122, 8'd10}: color_data = 12'hfd0;
			{8'd122, 8'd11}: color_data = 12'hfd0;
			{8'd122, 8'd12}: color_data = 12'hfc0;
			{8'd122, 8'd13}: color_data = 12'hfc0;
			{8'd122, 8'd14}: color_data = 12'hfc0;
			{8'd122, 8'd15}: color_data = 12'hfc0;
			{8'd122, 8'd16}: color_data = 12'hfc0;
			{8'd122, 8'd17}: color_data = 12'hfc0;
			{8'd122, 8'd18}: color_data = 12'hfd0;
			{8'd122, 8'd19}: color_data = 12'hfd0;
			{8'd122, 8'd20}: color_data = 12'hfd0;
			{8'd122, 8'd21}: color_data = 12'hfd0;
			{8'd122, 8'd22}: color_data = 12'hfd0;
			{8'd122, 8'd23}: color_data = 12'hfd0;
			{8'd122, 8'd24}: color_data = 12'hfd0;
			{8'd122, 8'd25}: color_data = 12'hfd0;
			{8'd122, 8'd26}: color_data = 12'hfd0;
			{8'd122, 8'd27}: color_data = 12'hfd0;
			{8'd122, 8'd28}: color_data = 12'hfc0;
			{8'd122, 8'd29}: color_data = 12'hfc0;
			{8'd122, 8'd30}: color_data = 12'hb90;
			{8'd122, 8'd31}: color_data = 12'h000;
			{8'd122, 8'd32}: color_data = 12'h000;
			{8'd122, 8'd33}: color_data = 12'h000;
			{8'd122, 8'd34}: color_data = 12'h000;
			{8'd122, 8'd35}: color_data = 12'h000;
			{8'd122, 8'd36}: color_data = 12'h08b;
			{8'd122, 8'd37}: color_data = 12'h09d;
			{8'd122, 8'd38}: color_data = 12'h09d;
			{8'd122, 8'd39}: color_data = 12'h09d;
			{8'd122, 8'd40}: color_data = 12'h09d;
			{8'd122, 8'd41}: color_data = 12'h09d;
			{8'd122, 8'd42}: color_data = 12'h09d;
			{8'd122, 8'd43}: color_data = 12'h09d;
			{8'd122, 8'd44}: color_data = 12'h09d;
			{8'd122, 8'd45}: color_data = 12'h09d;
			{8'd122, 8'd46}: color_data = 12'h09d;
			{8'd122, 8'd47}: color_data = 12'h09d;
			{8'd122, 8'd48}: color_data = 12'h09d;
			{8'd122, 8'd49}: color_data = 12'h09d;
			{8'd122, 8'd50}: color_data = 12'h0ae;
			{8'd122, 8'd51}: color_data = 12'h0ae;
			{8'd122, 8'd52}: color_data = 12'h09d;
			{8'd122, 8'd53}: color_data = 12'h09d;
			{8'd122, 8'd54}: color_data = 12'h08c;
			{8'd122, 8'd55}: color_data = 12'h07a;
			{8'd122, 8'd56}: color_data = 12'h058;
			{8'd122, 8'd57}: color_data = 12'h045;
			{8'd122, 8'd58}: color_data = 12'h023;
			{8'd122, 8'd59}: color_data = 12'h011;
			{8'd122, 8'd60}: color_data = 12'h000;
			{8'd122, 8'd61}: color_data = 12'h000;
			{8'd122, 8'd62}: color_data = 12'h000;
			{8'd122, 8'd63}: color_data = 12'h000;
			{8'd122, 8'd64}: color_data = 12'h000;
			{8'd122, 8'd65}: color_data = 12'h000;
			{8'd122, 8'd66}: color_data = 12'h000;
			{8'd122, 8'd67}: color_data = 12'h000;
			{8'd122, 8'd68}: color_data = 12'h000;
			{8'd122, 8'd69}: color_data = 12'h000;
			{8'd122, 8'd70}: color_data = 12'h000;
			{8'd122, 8'd71}: color_data = 12'h000;
			{8'd122, 8'd72}: color_data = 12'h000;
			{8'd122, 8'd73}: color_data = 12'h000;
			{8'd122, 8'd74}: color_data = 12'h000;
			{8'd122, 8'd100}: color_data = 12'he00;
			{8'd122, 8'd101}: color_data = 12'hf01;
			{8'd122, 8'd102}: color_data = 12'he00;
			{8'd122, 8'd103}: color_data = 12'he00;
			{8'd122, 8'd104}: color_data = 12'he00;
			{8'd122, 8'd105}: color_data = 12'he00;
			{8'd122, 8'd106}: color_data = 12'hc00;
			{8'd122, 8'd138}: color_data = 12'he00;
			{8'd122, 8'd139}: color_data = 12'he00;
			{8'd122, 8'd140}: color_data = 12'he00;
			{8'd122, 8'd141}: color_data = 12'he00;
			{8'd122, 8'd142}: color_data = 12'he00;
			{8'd122, 8'd143}: color_data = 12'he01;
			{8'd122, 8'd144}: color_data = 12'he00;
			{8'd123, 8'd2}: color_data = 12'h000;
			{8'd123, 8'd3}: color_data = 12'h000;
			{8'd123, 8'd4}: color_data = 12'h220;
			{8'd123, 8'd5}: color_data = 12'hfc0;
			{8'd123, 8'd6}: color_data = 12'hfd0;
			{8'd123, 8'd7}: color_data = 12'hfc0;
			{8'd123, 8'd8}: color_data = 12'hfc0;
			{8'd123, 8'd9}: color_data = 12'hfc0;
			{8'd123, 8'd10}: color_data = 12'hfc0;
			{8'd123, 8'd11}: color_data = 12'hfc0;
			{8'd123, 8'd12}: color_data = 12'hfc0;
			{8'd123, 8'd13}: color_data = 12'hfc0;
			{8'd123, 8'd14}: color_data = 12'hfc0;
			{8'd123, 8'd15}: color_data = 12'hfc0;
			{8'd123, 8'd16}: color_data = 12'hfc0;
			{8'd123, 8'd17}: color_data = 12'hfc0;
			{8'd123, 8'd18}: color_data = 12'hfc0;
			{8'd123, 8'd19}: color_data = 12'hfc0;
			{8'd123, 8'd20}: color_data = 12'hfc0;
			{8'd123, 8'd21}: color_data = 12'hfc0;
			{8'd123, 8'd22}: color_data = 12'hfc0;
			{8'd123, 8'd23}: color_data = 12'hfc0;
			{8'd123, 8'd24}: color_data = 12'hfc0;
			{8'd123, 8'd25}: color_data = 12'hfc0;
			{8'd123, 8'd26}: color_data = 12'hfc0;
			{8'd123, 8'd27}: color_data = 12'hfd0;
			{8'd123, 8'd28}: color_data = 12'hfd0;
			{8'd123, 8'd29}: color_data = 12'hfd0;
			{8'd123, 8'd30}: color_data = 12'hca0;
			{8'd123, 8'd31}: color_data = 12'h000;
			{8'd123, 8'd32}: color_data = 12'h000;
			{8'd123, 8'd33}: color_data = 12'h000;
			{8'd123, 8'd34}: color_data = 12'h000;
			{8'd123, 8'd35}: color_data = 12'h000;
			{8'd123, 8'd36}: color_data = 12'h069;
			{8'd123, 8'd37}: color_data = 12'h0ae;
			{8'd123, 8'd38}: color_data = 12'h09d;
			{8'd123, 8'd39}: color_data = 12'h09d;
			{8'd123, 8'd40}: color_data = 12'h09d;
			{8'd123, 8'd41}: color_data = 12'h09d;
			{8'd123, 8'd42}: color_data = 12'h09d;
			{8'd123, 8'd43}: color_data = 12'h09d;
			{8'd123, 8'd44}: color_data = 12'h0ae;
			{8'd123, 8'd45}: color_data = 12'h0ae;
			{8'd123, 8'd46}: color_data = 12'h0ae;
			{8'd123, 8'd47}: color_data = 12'h09d;
			{8'd123, 8'd48}: color_data = 12'h08c;
			{8'd123, 8'd49}: color_data = 12'h07a;
			{8'd123, 8'd50}: color_data = 12'h068;
			{8'd123, 8'd51}: color_data = 12'h046;
			{8'd123, 8'd52}: color_data = 12'h034;
			{8'd123, 8'd53}: color_data = 12'h012;
			{8'd123, 8'd54}: color_data = 12'h000;
			{8'd123, 8'd55}: color_data = 12'h000;
			{8'd123, 8'd56}: color_data = 12'h000;
			{8'd123, 8'd57}: color_data = 12'h000;
			{8'd123, 8'd58}: color_data = 12'h000;
			{8'd123, 8'd59}: color_data = 12'h000;
			{8'd123, 8'd60}: color_data = 12'h000;
			{8'd123, 8'd61}: color_data = 12'h000;
			{8'd123, 8'd62}: color_data = 12'h000;
			{8'd123, 8'd63}: color_data = 12'h000;
			{8'd123, 8'd64}: color_data = 12'h000;
			{8'd123, 8'd65}: color_data = 12'h000;
			{8'd123, 8'd66}: color_data = 12'h000;
			{8'd123, 8'd67}: color_data = 12'h000;
			{8'd123, 8'd68}: color_data = 12'h000;
			{8'd123, 8'd69}: color_data = 12'h000;
			{8'd123, 8'd70}: color_data = 12'h000;
			{8'd123, 8'd71}: color_data = 12'h000;
			{8'd123, 8'd72}: color_data = 12'h000;
			{8'd123, 8'd73}: color_data = 12'h000;
			{8'd123, 8'd100}: color_data = 12'he00;
			{8'd123, 8'd101}: color_data = 12'hf01;
			{8'd123, 8'd102}: color_data = 12'he00;
			{8'd123, 8'd103}: color_data = 12'he00;
			{8'd123, 8'd104}: color_data = 12'he00;
			{8'd123, 8'd105}: color_data = 12'he00;
			{8'd123, 8'd106}: color_data = 12'hc00;
			{8'd123, 8'd122}: color_data = 12'hf00;
			{8'd123, 8'd123}: color_data = 12'he00;
			{8'd123, 8'd124}: color_data = 12'he00;
			{8'd123, 8'd125}: color_data = 12'he01;
			{8'd123, 8'd126}: color_data = 12'he00;
			{8'd123, 8'd127}: color_data = 12'he00;
			{8'd123, 8'd128}: color_data = 12'hd01;
			{8'd123, 8'd138}: color_data = 12'he00;
			{8'd123, 8'd139}: color_data = 12'he00;
			{8'd123, 8'd140}: color_data = 12'he00;
			{8'd123, 8'd141}: color_data = 12'he00;
			{8'd123, 8'd142}: color_data = 12'he00;
			{8'd123, 8'd143}: color_data = 12'he01;
			{8'd123, 8'd144}: color_data = 12'he00;
			{8'd124, 8'd2}: color_data = 12'h000;
			{8'd124, 8'd3}: color_data = 12'h000;
			{8'd124, 8'd4}: color_data = 12'h430;
			{8'd124, 8'd5}: color_data = 12'hfd0;
			{8'd124, 8'd6}: color_data = 12'hfc0;
			{8'd124, 8'd7}: color_data = 12'hfc0;
			{8'd124, 8'd8}: color_data = 12'hfc0;
			{8'd124, 8'd9}: color_data = 12'hfc0;
			{8'd124, 8'd10}: color_data = 12'hfc0;
			{8'd124, 8'd11}: color_data = 12'hfc0;
			{8'd124, 8'd12}: color_data = 12'hfc0;
			{8'd124, 8'd13}: color_data = 12'hfc0;
			{8'd124, 8'd14}: color_data = 12'hfc0;
			{8'd124, 8'd15}: color_data = 12'hfc0;
			{8'd124, 8'd16}: color_data = 12'hfc0;
			{8'd124, 8'd17}: color_data = 12'hfc0;
			{8'd124, 8'd18}: color_data = 12'hfc0;
			{8'd124, 8'd19}: color_data = 12'hfc0;
			{8'd124, 8'd20}: color_data = 12'hfc0;
			{8'd124, 8'd21}: color_data = 12'hfc0;
			{8'd124, 8'd22}: color_data = 12'hfc0;
			{8'd124, 8'd23}: color_data = 12'hfc0;
			{8'd124, 8'd24}: color_data = 12'hfc0;
			{8'd124, 8'd25}: color_data = 12'hfc0;
			{8'd124, 8'd26}: color_data = 12'hfc0;
			{8'd124, 8'd27}: color_data = 12'hfc0;
			{8'd124, 8'd28}: color_data = 12'hfc0;
			{8'd124, 8'd29}: color_data = 12'hfd0;
			{8'd124, 8'd30}: color_data = 12'ha90;
			{8'd124, 8'd31}: color_data = 12'h000;
			{8'd124, 8'd32}: color_data = 12'h000;
			{8'd124, 8'd33}: color_data = 12'h000;
			{8'd124, 8'd34}: color_data = 12'h000;
			{8'd124, 8'd35}: color_data = 12'h000;
			{8'd124, 8'd36}: color_data = 12'h046;
			{8'd124, 8'd37}: color_data = 12'h0ae;
			{8'd124, 8'd38}: color_data = 12'h09d;
			{8'd124, 8'd39}: color_data = 12'h0ae;
			{8'd124, 8'd40}: color_data = 12'h0ae;
			{8'd124, 8'd41}: color_data = 12'h09d;
			{8'd124, 8'd42}: color_data = 12'h09c;
			{8'd124, 8'd43}: color_data = 12'h08b;
			{8'd124, 8'd44}: color_data = 12'h069;
			{8'd124, 8'd45}: color_data = 12'h057;
			{8'd124, 8'd46}: color_data = 12'h035;
			{8'd124, 8'd47}: color_data = 12'h022;
			{8'd124, 8'd48}: color_data = 12'h001;
			{8'd124, 8'd49}: color_data = 12'h000;
			{8'd124, 8'd50}: color_data = 12'h000;
			{8'd124, 8'd51}: color_data = 12'h000;
			{8'd124, 8'd52}: color_data = 12'h000;
			{8'd124, 8'd53}: color_data = 12'h000;
			{8'd124, 8'd54}: color_data = 12'h000;
			{8'd124, 8'd55}: color_data = 12'h000;
			{8'd124, 8'd56}: color_data = 12'h000;
			{8'd124, 8'd57}: color_data = 12'h000;
			{8'd124, 8'd58}: color_data = 12'h000;
			{8'd124, 8'd59}: color_data = 12'h000;
			{8'd124, 8'd60}: color_data = 12'h000;
			{8'd124, 8'd61}: color_data = 12'h000;
			{8'd124, 8'd62}: color_data = 12'h000;
			{8'd124, 8'd63}: color_data = 12'h000;
			{8'd124, 8'd64}: color_data = 12'h000;
			{8'd124, 8'd65}: color_data = 12'h000;
			{8'd124, 8'd66}: color_data = 12'h000;
			{8'd124, 8'd67}: color_data = 12'h000;
			{8'd124, 8'd100}: color_data = 12'he00;
			{8'd124, 8'd101}: color_data = 12'hf01;
			{8'd124, 8'd102}: color_data = 12'he00;
			{8'd124, 8'd103}: color_data = 12'he00;
			{8'd124, 8'd104}: color_data = 12'he00;
			{8'd124, 8'd105}: color_data = 12'he00;
			{8'd124, 8'd106}: color_data = 12'hc00;
			{8'd124, 8'd121}: color_data = 12'he00;
			{8'd124, 8'd122}: color_data = 12'he00;
			{8'd124, 8'd123}: color_data = 12'he00;
			{8'd124, 8'd124}: color_data = 12'he00;
			{8'd124, 8'd125}: color_data = 12'he00;
			{8'd124, 8'd126}: color_data = 12'he00;
			{8'd124, 8'd127}: color_data = 12'he00;
			{8'd124, 8'd128}: color_data = 12'he00;
			{8'd124, 8'd129}: color_data = 12'he00;
			{8'd124, 8'd130}: color_data = 12'he00;
			{8'd124, 8'd138}: color_data = 12'he00;
			{8'd124, 8'd139}: color_data = 12'he00;
			{8'd124, 8'd140}: color_data = 12'he00;
			{8'd124, 8'd141}: color_data = 12'he00;
			{8'd124, 8'd142}: color_data = 12'he00;
			{8'd124, 8'd143}: color_data = 12'he01;
			{8'd124, 8'd144}: color_data = 12'he00;
			{8'd125, 8'd2}: color_data = 12'h000;
			{8'd125, 8'd3}: color_data = 12'h000;
			{8'd125, 8'd4}: color_data = 12'h650;
			{8'd125, 8'd5}: color_data = 12'hfd0;
			{8'd125, 8'd6}: color_data = 12'hfc0;
			{8'd125, 8'd7}: color_data = 12'hfc0;
			{8'd125, 8'd8}: color_data = 12'hfc0;
			{8'd125, 8'd9}: color_data = 12'hfc0;
			{8'd125, 8'd10}: color_data = 12'hfc0;
			{8'd125, 8'd11}: color_data = 12'hfc0;
			{8'd125, 8'd12}: color_data = 12'hfc0;
			{8'd125, 8'd13}: color_data = 12'hfc0;
			{8'd125, 8'd14}: color_data = 12'hfc0;
			{8'd125, 8'd15}: color_data = 12'hfc0;
			{8'd125, 8'd16}: color_data = 12'hfc0;
			{8'd125, 8'd17}: color_data = 12'hfc0;
			{8'd125, 8'd18}: color_data = 12'hfc0;
			{8'd125, 8'd19}: color_data = 12'hfc0;
			{8'd125, 8'd20}: color_data = 12'hfc0;
			{8'd125, 8'd21}: color_data = 12'hfc0;
			{8'd125, 8'd22}: color_data = 12'hfc0;
			{8'd125, 8'd23}: color_data = 12'hfc0;
			{8'd125, 8'd24}: color_data = 12'hfc0;
			{8'd125, 8'd25}: color_data = 12'hfc0;
			{8'd125, 8'd26}: color_data = 12'hfc0;
			{8'd125, 8'd27}: color_data = 12'hfc0;
			{8'd125, 8'd28}: color_data = 12'hfc0;
			{8'd125, 8'd29}: color_data = 12'hfd0;
			{8'd125, 8'd30}: color_data = 12'h980;
			{8'd125, 8'd31}: color_data = 12'h000;
			{8'd125, 8'd32}: color_data = 12'h000;
			{8'd125, 8'd33}: color_data = 12'h000;
			{8'd125, 8'd34}: color_data = 12'h000;
			{8'd125, 8'd35}: color_data = 12'h000;
			{8'd125, 8'd36}: color_data = 12'h022;
			{8'd125, 8'd37}: color_data = 12'h08b;
			{8'd125, 8'd38}: color_data = 12'h07a;
			{8'd125, 8'd39}: color_data = 12'h058;
			{8'd125, 8'd40}: color_data = 12'h045;
			{8'd125, 8'd41}: color_data = 12'h023;
			{8'd125, 8'd42}: color_data = 12'h011;
			{8'd125, 8'd43}: color_data = 12'h000;
			{8'd125, 8'd44}: color_data = 12'h000;
			{8'd125, 8'd45}: color_data = 12'h000;
			{8'd125, 8'd46}: color_data = 12'h000;
			{8'd125, 8'd47}: color_data = 12'h000;
			{8'd125, 8'd48}: color_data = 12'h000;
			{8'd125, 8'd49}: color_data = 12'h000;
			{8'd125, 8'd50}: color_data = 12'h000;
			{8'd125, 8'd51}: color_data = 12'h000;
			{8'd125, 8'd52}: color_data = 12'h000;
			{8'd125, 8'd53}: color_data = 12'h020;
			{8'd125, 8'd54}: color_data = 12'h141;
			{8'd125, 8'd55}: color_data = 12'h141;
			{8'd125, 8'd56}: color_data = 12'h010;
			{8'd125, 8'd57}: color_data = 12'h000;
			{8'd125, 8'd58}: color_data = 12'h000;
			{8'd125, 8'd59}: color_data = 12'h000;
			{8'd125, 8'd60}: color_data = 12'h000;
			{8'd125, 8'd61}: color_data = 12'h000;
			{8'd125, 8'd62}: color_data = 12'h000;
			{8'd125, 8'd63}: color_data = 12'h000;
			{8'd125, 8'd64}: color_data = 12'h000;
			{8'd125, 8'd65}: color_data = 12'h000;
			{8'd125, 8'd66}: color_data = 12'h000;
			{8'd125, 8'd67}: color_data = 12'h000;
			{8'd125, 8'd68}: color_data = 12'h000;
			{8'd125, 8'd69}: color_data = 12'h000;
			{8'd125, 8'd100}: color_data = 12'he00;
			{8'd125, 8'd101}: color_data = 12'hf01;
			{8'd125, 8'd102}: color_data = 12'he00;
			{8'd125, 8'd103}: color_data = 12'he00;
			{8'd125, 8'd104}: color_data = 12'he00;
			{8'd125, 8'd105}: color_data = 12'he00;
			{8'd125, 8'd106}: color_data = 12'hc00;
			{8'd125, 8'd119}: color_data = 12'hc00;
			{8'd125, 8'd120}: color_data = 12'he00;
			{8'd125, 8'd121}: color_data = 12'he00;
			{8'd125, 8'd122}: color_data = 12'he00;
			{8'd125, 8'd123}: color_data = 12'he00;
			{8'd125, 8'd124}: color_data = 12'he00;
			{8'd125, 8'd125}: color_data = 12'he00;
			{8'd125, 8'd126}: color_data = 12'he00;
			{8'd125, 8'd127}: color_data = 12'he00;
			{8'd125, 8'd128}: color_data = 12'he00;
			{8'd125, 8'd129}: color_data = 12'hf01;
			{8'd125, 8'd130}: color_data = 12'he00;
			{8'd125, 8'd131}: color_data = 12'he00;
			{8'd125, 8'd138}: color_data = 12'he00;
			{8'd125, 8'd139}: color_data = 12'he00;
			{8'd125, 8'd140}: color_data = 12'he00;
			{8'd125, 8'd141}: color_data = 12'he00;
			{8'd125, 8'd142}: color_data = 12'he00;
			{8'd125, 8'd143}: color_data = 12'he01;
			{8'd125, 8'd144}: color_data = 12'he00;
			{8'd126, 8'd1}: color_data = 12'h000;
			{8'd126, 8'd2}: color_data = 12'h000;
			{8'd126, 8'd3}: color_data = 12'h000;
			{8'd126, 8'd4}: color_data = 12'h970;
			{8'd126, 8'd5}: color_data = 12'hfd0;
			{8'd126, 8'd6}: color_data = 12'hfc0;
			{8'd126, 8'd7}: color_data = 12'hfc0;
			{8'd126, 8'd8}: color_data = 12'hfc0;
			{8'd126, 8'd9}: color_data = 12'hfc0;
			{8'd126, 8'd10}: color_data = 12'hfc0;
			{8'd126, 8'd11}: color_data = 12'hfc0;
			{8'd126, 8'd12}: color_data = 12'hfc0;
			{8'd126, 8'd13}: color_data = 12'hfc0;
			{8'd126, 8'd14}: color_data = 12'hfc0;
			{8'd126, 8'd15}: color_data = 12'hfc0;
			{8'd126, 8'd16}: color_data = 12'hfc0;
			{8'd126, 8'd17}: color_data = 12'hfc0;
			{8'd126, 8'd18}: color_data = 12'hfc0;
			{8'd126, 8'd19}: color_data = 12'hfc0;
			{8'd126, 8'd20}: color_data = 12'hfc0;
			{8'd126, 8'd21}: color_data = 12'hfc0;
			{8'd126, 8'd22}: color_data = 12'hfc0;
			{8'd126, 8'd23}: color_data = 12'hfc0;
			{8'd126, 8'd24}: color_data = 12'hfc0;
			{8'd126, 8'd25}: color_data = 12'hfc0;
			{8'd126, 8'd26}: color_data = 12'hfc0;
			{8'd126, 8'd27}: color_data = 12'hfc0;
			{8'd126, 8'd28}: color_data = 12'hfc0;
			{8'd126, 8'd29}: color_data = 12'hfd0;
			{8'd126, 8'd30}: color_data = 12'h860;
			{8'd126, 8'd31}: color_data = 12'h000;
			{8'd126, 8'd32}: color_data = 12'h000;
			{8'd126, 8'd33}: color_data = 12'h000;
			{8'd126, 8'd34}: color_data = 12'h000;
			{8'd126, 8'd35}: color_data = 12'h000;
			{8'd126, 8'd36}: color_data = 12'h000;
			{8'd126, 8'd37}: color_data = 12'h000;
			{8'd126, 8'd38}: color_data = 12'h000;
			{8'd126, 8'd39}: color_data = 12'h000;
			{8'd126, 8'd40}: color_data = 12'h000;
			{8'd126, 8'd41}: color_data = 12'h000;
			{8'd126, 8'd42}: color_data = 12'h000;
			{8'd126, 8'd43}: color_data = 12'h000;
			{8'd126, 8'd44}: color_data = 12'h000;
			{8'd126, 8'd45}: color_data = 12'h000;
			{8'd126, 8'd46}: color_data = 12'h000;
			{8'd126, 8'd47}: color_data = 12'h010;
			{8'd126, 8'd48}: color_data = 12'h131;
			{8'd126, 8'd49}: color_data = 12'h151;
			{8'd126, 8'd50}: color_data = 12'h262;
			{8'd126, 8'd51}: color_data = 12'h382;
			{8'd126, 8'd52}: color_data = 12'h3a3;
			{8'd126, 8'd53}: color_data = 12'h4a3;
			{8'd126, 8'd54}: color_data = 12'h4b3;
			{8'd126, 8'd55}: color_data = 12'h4b3;
			{8'd126, 8'd56}: color_data = 12'h4a3;
			{8'd126, 8'd57}: color_data = 12'h382;
			{8'd126, 8'd58}: color_data = 12'h141;
			{8'd126, 8'd59}: color_data = 12'h010;
			{8'd126, 8'd60}: color_data = 12'h000;
			{8'd126, 8'd61}: color_data = 12'h000;
			{8'd126, 8'd62}: color_data = 12'h000;
			{8'd126, 8'd63}: color_data = 12'h000;
			{8'd126, 8'd64}: color_data = 12'h000;
			{8'd126, 8'd65}: color_data = 12'h000;
			{8'd126, 8'd66}: color_data = 12'h000;
			{8'd126, 8'd67}: color_data = 12'h000;
			{8'd126, 8'd68}: color_data = 12'h000;
			{8'd126, 8'd69}: color_data = 12'h000;
			{8'd126, 8'd70}: color_data = 12'h000;
			{8'd126, 8'd71}: color_data = 12'h000;
			{8'd126, 8'd100}: color_data = 12'he00;
			{8'd126, 8'd101}: color_data = 12'hf01;
			{8'd126, 8'd102}: color_data = 12'he00;
			{8'd126, 8'd103}: color_data = 12'he00;
			{8'd126, 8'd104}: color_data = 12'he00;
			{8'd126, 8'd105}: color_data = 12'he00;
			{8'd126, 8'd106}: color_data = 12'hc00;
			{8'd126, 8'd119}: color_data = 12'he00;
			{8'd126, 8'd120}: color_data = 12'hf01;
			{8'd126, 8'd121}: color_data = 12'he00;
			{8'd126, 8'd122}: color_data = 12'he00;
			{8'd126, 8'd123}: color_data = 12'he00;
			{8'd126, 8'd124}: color_data = 12'he00;
			{8'd126, 8'd125}: color_data = 12'he00;
			{8'd126, 8'd126}: color_data = 12'he00;
			{8'd126, 8'd127}: color_data = 12'he00;
			{8'd126, 8'd128}: color_data = 12'he00;
			{8'd126, 8'd129}: color_data = 12'he00;
			{8'd126, 8'd130}: color_data = 12'he01;
			{8'd126, 8'd131}: color_data = 12'he00;
			{8'd126, 8'd132}: color_data = 12'he00;
			{8'd126, 8'd138}: color_data = 12'he00;
			{8'd126, 8'd139}: color_data = 12'he00;
			{8'd126, 8'd140}: color_data = 12'he00;
			{8'd126, 8'd141}: color_data = 12'he00;
			{8'd126, 8'd142}: color_data = 12'he00;
			{8'd126, 8'd143}: color_data = 12'he01;
			{8'd126, 8'd144}: color_data = 12'he00;
			{8'd127, 8'd1}: color_data = 12'h000;
			{8'd127, 8'd2}: color_data = 12'h000;
			{8'd127, 8'd3}: color_data = 12'h000;
			{8'd127, 8'd4}: color_data = 12'hb90;
			{8'd127, 8'd5}: color_data = 12'hfd0;
			{8'd127, 8'd6}: color_data = 12'hfc0;
			{8'd127, 8'd7}: color_data = 12'hfc0;
			{8'd127, 8'd8}: color_data = 12'hfc0;
			{8'd127, 8'd9}: color_data = 12'hfd0;
			{8'd127, 8'd10}: color_data = 12'hfd0;
			{8'd127, 8'd11}: color_data = 12'hfd0;
			{8'd127, 8'd12}: color_data = 12'hfd0;
			{8'd127, 8'd13}: color_data = 12'hfd0;
			{8'd127, 8'd14}: color_data = 12'hfd0;
			{8'd127, 8'd15}: color_data = 12'hfd0;
			{8'd127, 8'd16}: color_data = 12'hfd0;
			{8'd127, 8'd17}: color_data = 12'hfd0;
			{8'd127, 8'd18}: color_data = 12'hfd0;
			{8'd127, 8'd19}: color_data = 12'hfc0;
			{8'd127, 8'd20}: color_data = 12'hfc0;
			{8'd127, 8'd21}: color_data = 12'hfd0;
			{8'd127, 8'd22}: color_data = 12'hfd0;
			{8'd127, 8'd23}: color_data = 12'hfd0;
			{8'd127, 8'd24}: color_data = 12'hfd0;
			{8'd127, 8'd25}: color_data = 12'hfd0;
			{8'd127, 8'd26}: color_data = 12'hfd0;
			{8'd127, 8'd27}: color_data = 12'hfd0;
			{8'd127, 8'd28}: color_data = 12'hfd0;
			{8'd127, 8'd29}: color_data = 12'hfd0;
			{8'd127, 8'd30}: color_data = 12'h650;
			{8'd127, 8'd31}: color_data = 12'h000;
			{8'd127, 8'd32}: color_data = 12'h000;
			{8'd127, 8'd33}: color_data = 12'h000;
			{8'd127, 8'd34}: color_data = 12'h000;
			{8'd127, 8'd35}: color_data = 12'h000;
			{8'd127, 8'd36}: color_data = 12'h000;
			{8'd127, 8'd37}: color_data = 12'h000;
			{8'd127, 8'd38}: color_data = 12'h000;
			{8'd127, 8'd39}: color_data = 12'h000;
			{8'd127, 8'd40}: color_data = 12'h000;
			{8'd127, 8'd41}: color_data = 12'h000;
			{8'd127, 8'd42}: color_data = 12'h000;
			{8'd127, 8'd43}: color_data = 12'h000;
			{8'd127, 8'd44}: color_data = 12'h251;
			{8'd127, 8'd45}: color_data = 12'h382;
			{8'd127, 8'd46}: color_data = 12'h392;
			{8'd127, 8'd47}: color_data = 12'h4a3;
			{8'd127, 8'd48}: color_data = 12'h4b3;
			{8'd127, 8'd49}: color_data = 12'h4b3;
			{8'd127, 8'd50}: color_data = 12'h4b3;
			{8'd127, 8'd51}: color_data = 12'h4b3;
			{8'd127, 8'd52}: color_data = 12'h4b3;
			{8'd127, 8'd53}: color_data = 12'h4b3;
			{8'd127, 8'd54}: color_data = 12'h4a3;
			{8'd127, 8'd55}: color_data = 12'h4a3;
			{8'd127, 8'd56}: color_data = 12'h4b3;
			{8'd127, 8'd57}: color_data = 12'h4b3;
			{8'd127, 8'd58}: color_data = 12'h4b3;
			{8'd127, 8'd59}: color_data = 12'h4a3;
			{8'd127, 8'd60}: color_data = 12'h372;
			{8'd127, 8'd61}: color_data = 12'h141;
			{8'd127, 8'd62}: color_data = 12'h010;
			{8'd127, 8'd63}: color_data = 12'h000;
			{8'd127, 8'd64}: color_data = 12'h000;
			{8'd127, 8'd65}: color_data = 12'h000;
			{8'd127, 8'd66}: color_data = 12'h000;
			{8'd127, 8'd67}: color_data = 12'h000;
			{8'd127, 8'd68}: color_data = 12'h000;
			{8'd127, 8'd69}: color_data = 12'h000;
			{8'd127, 8'd70}: color_data = 12'h000;
			{8'd127, 8'd71}: color_data = 12'h000;
			{8'd127, 8'd100}: color_data = 12'he00;
			{8'd127, 8'd101}: color_data = 12'hf01;
			{8'd127, 8'd102}: color_data = 12'he00;
			{8'd127, 8'd103}: color_data = 12'he00;
			{8'd127, 8'd104}: color_data = 12'he00;
			{8'd127, 8'd105}: color_data = 12'he00;
			{8'd127, 8'd106}: color_data = 12'hc00;
			{8'd127, 8'd118}: color_data = 12'he00;
			{8'd127, 8'd119}: color_data = 12'he00;
			{8'd127, 8'd120}: color_data = 12'he00;
			{8'd127, 8'd121}: color_data = 12'he00;
			{8'd127, 8'd122}: color_data = 12'he00;
			{8'd127, 8'd123}: color_data = 12'he00;
			{8'd127, 8'd124}: color_data = 12'he00;
			{8'd127, 8'd125}: color_data = 12'he00;
			{8'd127, 8'd126}: color_data = 12'he00;
			{8'd127, 8'd127}: color_data = 12'he00;
			{8'd127, 8'd128}: color_data = 12'he00;
			{8'd127, 8'd129}: color_data = 12'he00;
			{8'd127, 8'd130}: color_data = 12'he00;
			{8'd127, 8'd131}: color_data = 12'hf01;
			{8'd127, 8'd132}: color_data = 12'he00;
			{8'd127, 8'd138}: color_data = 12'he00;
			{8'd127, 8'd139}: color_data = 12'he00;
			{8'd127, 8'd140}: color_data = 12'he00;
			{8'd127, 8'd141}: color_data = 12'he00;
			{8'd127, 8'd142}: color_data = 12'he00;
			{8'd127, 8'd143}: color_data = 12'he01;
			{8'd127, 8'd144}: color_data = 12'he00;
			{8'd128, 8'd1}: color_data = 12'h000;
			{8'd128, 8'd2}: color_data = 12'h000;
			{8'd128, 8'd3}: color_data = 12'h000;
			{8'd128, 8'd4}: color_data = 12'hda0;
			{8'd128, 8'd5}: color_data = 12'hfd0;
			{8'd128, 8'd6}: color_data = 12'hfc0;
			{8'd128, 8'd7}: color_data = 12'hfc0;
			{8'd128, 8'd8}: color_data = 12'hfd0;
			{8'd128, 8'd9}: color_data = 12'heb0;
			{8'd128, 8'd10}: color_data = 12'h750;
			{8'd128, 8'd11}: color_data = 12'h750;
			{8'd128, 8'd12}: color_data = 12'h760;
			{8'd128, 8'd13}: color_data = 12'h860;
			{8'd128, 8'd14}: color_data = 12'h870;
			{8'd128, 8'd15}: color_data = 12'h970;
			{8'd128, 8'd16}: color_data = 12'h970;
			{8'd128, 8'd17}: color_data = 12'ha80;
			{8'd128, 8'd18}: color_data = 12'hec0;
			{8'd128, 8'd19}: color_data = 12'hfd0;
			{8'd128, 8'd20}: color_data = 12'hfd0;
			{8'd128, 8'd21}: color_data = 12'hfc0;
			{8'd128, 8'd22}: color_data = 12'hc90;
			{8'd128, 8'd23}: color_data = 12'hca0;
			{8'd128, 8'd24}: color_data = 12'hda0;
			{8'd128, 8'd25}: color_data = 12'hda0;
			{8'd128, 8'd26}: color_data = 12'hdb0;
			{8'd128, 8'd27}: color_data = 12'heb0;
			{8'd128, 8'd28}: color_data = 12'heb0;
			{8'd128, 8'd29}: color_data = 12'hec0;
			{8'd128, 8'd30}: color_data = 12'h540;
			{8'd128, 8'd31}: color_data = 12'h000;
			{8'd128, 8'd32}: color_data = 12'h000;
			{8'd128, 8'd33}: color_data = 12'h000;
			{8'd128, 8'd34}: color_data = 12'h000;
			{8'd128, 8'd35}: color_data = 12'h000;
			{8'd128, 8'd36}: color_data = 12'h000;
			{8'd128, 8'd37}: color_data = 12'h000;
			{8'd128, 8'd38}: color_data = 12'h000;
			{8'd128, 8'd39}: color_data = 12'h000;
			{8'd128, 8'd40}: color_data = 12'h000;
			{8'd128, 8'd41}: color_data = 12'h000;
			{8'd128, 8'd42}: color_data = 12'h010;
			{8'd128, 8'd43}: color_data = 12'h382;
			{8'd128, 8'd44}: color_data = 12'h4b3;
			{8'd128, 8'd45}: color_data = 12'h4b3;
			{8'd128, 8'd46}: color_data = 12'h4b3;
			{8'd128, 8'd47}: color_data = 12'h4b3;
			{8'd128, 8'd48}: color_data = 12'h4a3;
			{8'd128, 8'd49}: color_data = 12'h4a3;
			{8'd128, 8'd50}: color_data = 12'h4a3;
			{8'd128, 8'd51}: color_data = 12'h4a3;
			{8'd128, 8'd52}: color_data = 12'h4a3;
			{8'd128, 8'd53}: color_data = 12'h4a3;
			{8'd128, 8'd54}: color_data = 12'h4a3;
			{8'd128, 8'd55}: color_data = 12'h4a3;
			{8'd128, 8'd56}: color_data = 12'h4a3;
			{8'd128, 8'd57}: color_data = 12'h4a3;
			{8'd128, 8'd58}: color_data = 12'h4a3;
			{8'd128, 8'd59}: color_data = 12'h4b3;
			{8'd128, 8'd60}: color_data = 12'h4b3;
			{8'd128, 8'd61}: color_data = 12'h4b3;
			{8'd128, 8'd62}: color_data = 12'h3a3;
			{8'd128, 8'd63}: color_data = 12'h272;
			{8'd128, 8'd64}: color_data = 12'h131;
			{8'd128, 8'd65}: color_data = 12'h000;
			{8'd128, 8'd66}: color_data = 12'h000;
			{8'd128, 8'd67}: color_data = 12'h000;
			{8'd128, 8'd68}: color_data = 12'h000;
			{8'd128, 8'd69}: color_data = 12'h000;
			{8'd128, 8'd70}: color_data = 12'h000;
			{8'd128, 8'd71}: color_data = 12'h000;
			{8'd128, 8'd72}: color_data = 12'h000;
			{8'd128, 8'd100}: color_data = 12'he00;
			{8'd128, 8'd101}: color_data = 12'hf01;
			{8'd128, 8'd102}: color_data = 12'he00;
			{8'd128, 8'd103}: color_data = 12'he00;
			{8'd128, 8'd104}: color_data = 12'he00;
			{8'd128, 8'd105}: color_data = 12'he00;
			{8'd128, 8'd106}: color_data = 12'hc00;
			{8'd128, 8'd118}: color_data = 12'he00;
			{8'd128, 8'd119}: color_data = 12'he01;
			{8'd128, 8'd120}: color_data = 12'he00;
			{8'd128, 8'd121}: color_data = 12'he00;
			{8'd128, 8'd122}: color_data = 12'he00;
			{8'd128, 8'd123}: color_data = 12'he00;
			{8'd128, 8'd124}: color_data = 12'he00;
			{8'd128, 8'd125}: color_data = 12'he01;
			{8'd128, 8'd126}: color_data = 12'he01;
			{8'd128, 8'd127}: color_data = 12'he00;
			{8'd128, 8'd128}: color_data = 12'he00;
			{8'd128, 8'd129}: color_data = 12'he00;
			{8'd128, 8'd130}: color_data = 12'he00;
			{8'd128, 8'd131}: color_data = 12'he00;
			{8'd128, 8'd132}: color_data = 12'he00;
			{8'd128, 8'd133}: color_data = 12'he00;
			{8'd128, 8'd138}: color_data = 12'he00;
			{8'd128, 8'd139}: color_data = 12'he00;
			{8'd128, 8'd140}: color_data = 12'he00;
			{8'd128, 8'd141}: color_data = 12'he00;
			{8'd128, 8'd142}: color_data = 12'he00;
			{8'd128, 8'd143}: color_data = 12'he01;
			{8'd128, 8'd144}: color_data = 12'he00;
			{8'd129, 8'd1}: color_data = 12'h000;
			{8'd129, 8'd2}: color_data = 12'h000;
			{8'd129, 8'd3}: color_data = 12'h110;
			{8'd129, 8'd4}: color_data = 12'hec0;
			{8'd129, 8'd5}: color_data = 12'hfd0;
			{8'd129, 8'd6}: color_data = 12'hfc0;
			{8'd129, 8'd7}: color_data = 12'hfc0;
			{8'd129, 8'd8}: color_data = 12'hfd0;
			{8'd129, 8'd9}: color_data = 12'hfc0;
			{8'd129, 8'd10}: color_data = 12'h220;
			{8'd129, 8'd11}: color_data = 12'h000;
			{8'd129, 8'd12}: color_data = 12'h000;
			{8'd129, 8'd13}: color_data = 12'h000;
			{8'd129, 8'd14}: color_data = 12'h000;
			{8'd129, 8'd15}: color_data = 12'h000;
			{8'd129, 8'd16}: color_data = 12'h000;
			{8'd129, 8'd17}: color_data = 12'h110;
			{8'd129, 8'd18}: color_data = 12'heb0;
			{8'd129, 8'd19}: color_data = 12'hfd0;
			{8'd129, 8'd20}: color_data = 12'hfd0;
			{8'd129, 8'd21}: color_data = 12'hfc0;
			{8'd129, 8'd22}: color_data = 12'h870;
			{8'd129, 8'd23}: color_data = 12'h100;
			{8'd129, 8'd24}: color_data = 12'h000;
			{8'd129, 8'd25}: color_data = 12'h000;
			{8'd129, 8'd26}: color_data = 12'h000;
			{8'd129, 8'd27}: color_data = 12'h000;
			{8'd129, 8'd28}: color_data = 12'h100;
			{8'd129, 8'd29}: color_data = 12'h110;
			{8'd129, 8'd30}: color_data = 12'h000;
			{8'd129, 8'd31}: color_data = 12'h000;
			{8'd129, 8'd32}: color_data = 12'h000;
			{8'd129, 8'd33}: color_data = 12'h000;
			{8'd129, 8'd34}: color_data = 12'h000;
			{8'd129, 8'd35}: color_data = 12'h000;
			{8'd129, 8'd36}: color_data = 12'h000;
			{8'd129, 8'd37}: color_data = 12'h000;
			{8'd129, 8'd38}: color_data = 12'h000;
			{8'd129, 8'd39}: color_data = 12'h000;
			{8'd129, 8'd40}: color_data = 12'h000;
			{8'd129, 8'd41}: color_data = 12'h130;
			{8'd129, 8'd42}: color_data = 12'h393;
			{8'd129, 8'd43}: color_data = 12'h4b3;
			{8'd129, 8'd44}: color_data = 12'h4a3;
			{8'd129, 8'd45}: color_data = 12'h4a3;
			{8'd129, 8'd46}: color_data = 12'h4a3;
			{8'd129, 8'd47}: color_data = 12'h4a3;
			{8'd129, 8'd48}: color_data = 12'h4a3;
			{8'd129, 8'd49}: color_data = 12'h4a3;
			{8'd129, 8'd50}: color_data = 12'h4a3;
			{8'd129, 8'd51}: color_data = 12'h4a3;
			{8'd129, 8'd52}: color_data = 12'h4a3;
			{8'd129, 8'd53}: color_data = 12'h4a3;
			{8'd129, 8'd54}: color_data = 12'h4a3;
			{8'd129, 8'd55}: color_data = 12'h4a3;
			{8'd129, 8'd56}: color_data = 12'h4a3;
			{8'd129, 8'd57}: color_data = 12'h4a3;
			{8'd129, 8'd58}: color_data = 12'h4a3;
			{8'd129, 8'd59}: color_data = 12'h4a3;
			{8'd129, 8'd60}: color_data = 12'h4a3;
			{8'd129, 8'd61}: color_data = 12'h4a3;
			{8'd129, 8'd62}: color_data = 12'h4b3;
			{8'd129, 8'd63}: color_data = 12'h4b3;
			{8'd129, 8'd64}: color_data = 12'h4b3;
			{8'd129, 8'd65}: color_data = 12'h141;
			{8'd129, 8'd66}: color_data = 12'h000;
			{8'd129, 8'd67}: color_data = 12'h000;
			{8'd129, 8'd68}: color_data = 12'h000;
			{8'd129, 8'd69}: color_data = 12'h000;
			{8'd129, 8'd70}: color_data = 12'h000;
			{8'd129, 8'd71}: color_data = 12'h000;
			{8'd129, 8'd72}: color_data = 12'h000;
			{8'd129, 8'd100}: color_data = 12'he00;
			{8'd129, 8'd101}: color_data = 12'hf01;
			{8'd129, 8'd102}: color_data = 12'he00;
			{8'd129, 8'd103}: color_data = 12'he00;
			{8'd129, 8'd104}: color_data = 12'he00;
			{8'd129, 8'd105}: color_data = 12'he00;
			{8'd129, 8'd106}: color_data = 12'hc00;
			{8'd129, 8'd117}: color_data = 12'he00;
			{8'd129, 8'd118}: color_data = 12'he00;
			{8'd129, 8'd119}: color_data = 12'he00;
			{8'd129, 8'd120}: color_data = 12'he00;
			{8'd129, 8'd121}: color_data = 12'he00;
			{8'd129, 8'd122}: color_data = 12'he00;
			{8'd129, 8'd123}: color_data = 12'he00;
			{8'd129, 8'd124}: color_data = 12'he00;
			{8'd129, 8'd125}: color_data = 12'he00;
			{8'd129, 8'd126}: color_data = 12'he00;
			{8'd129, 8'd127}: color_data = 12'he00;
			{8'd129, 8'd128}: color_data = 12'he00;
			{8'd129, 8'd129}: color_data = 12'he00;
			{8'd129, 8'd130}: color_data = 12'he00;
			{8'd129, 8'd131}: color_data = 12'he00;
			{8'd129, 8'd132}: color_data = 12'hf01;
			{8'd129, 8'd133}: color_data = 12'he00;
			{8'd129, 8'd138}: color_data = 12'he00;
			{8'd129, 8'd139}: color_data = 12'he00;
			{8'd129, 8'd140}: color_data = 12'he00;
			{8'd129, 8'd141}: color_data = 12'he00;
			{8'd129, 8'd142}: color_data = 12'he00;
			{8'd129, 8'd143}: color_data = 12'he01;
			{8'd129, 8'd144}: color_data = 12'he00;
			{8'd130, 8'd1}: color_data = 12'h000;
			{8'd130, 8'd2}: color_data = 12'h000;
			{8'd130, 8'd3}: color_data = 12'h320;
			{8'd130, 8'd4}: color_data = 12'hfc0;
			{8'd130, 8'd5}: color_data = 12'hfd0;
			{8'd130, 8'd6}: color_data = 12'hfc0;
			{8'd130, 8'd7}: color_data = 12'hfc0;
			{8'd130, 8'd8}: color_data = 12'hfc0;
			{8'd130, 8'd9}: color_data = 12'hfd0;
			{8'd130, 8'd10}: color_data = 12'h860;
			{8'd130, 8'd11}: color_data = 12'h000;
			{8'd130, 8'd12}: color_data = 12'h000;
			{8'd130, 8'd13}: color_data = 12'h000;
			{8'd130, 8'd14}: color_data = 12'h000;
			{8'd130, 8'd15}: color_data = 12'h000;
			{8'd130, 8'd16}: color_data = 12'h000;
			{8'd130, 8'd17}: color_data = 12'h320;
			{8'd130, 8'd18}: color_data = 12'hfc0;
			{8'd130, 8'd19}: color_data = 12'hfd0;
			{8'd130, 8'd20}: color_data = 12'hfc0;
			{8'd130, 8'd21}: color_data = 12'hfd0;
			{8'd130, 8'd22}: color_data = 12'hfd0;
			{8'd130, 8'd23}: color_data = 12'hda0;
			{8'd130, 8'd24}: color_data = 12'h430;
			{8'd130, 8'd25}: color_data = 12'h000;
			{8'd130, 8'd26}: color_data = 12'h000;
			{8'd130, 8'd27}: color_data = 12'h000;
			{8'd130, 8'd28}: color_data = 12'h000;
			{8'd130, 8'd29}: color_data = 12'h000;
			{8'd130, 8'd30}: color_data = 12'h000;
			{8'd130, 8'd31}: color_data = 12'h000;
			{8'd130, 8'd32}: color_data = 12'h000;
			{8'd130, 8'd33}: color_data = 12'h000;
			{8'd130, 8'd34}: color_data = 12'h000;
			{8'd130, 8'd35}: color_data = 12'h000;
			{8'd130, 8'd36}: color_data = 12'h000;
			{8'd130, 8'd37}: color_data = 12'h000;
			{8'd130, 8'd38}: color_data = 12'h000;
			{8'd130, 8'd39}: color_data = 12'h000;
			{8'd130, 8'd40}: color_data = 12'h251;
			{8'd130, 8'd41}: color_data = 12'h4a3;
			{8'd130, 8'd42}: color_data = 12'h4b3;
			{8'd130, 8'd43}: color_data = 12'h4a3;
			{8'd130, 8'd44}: color_data = 12'h4a3;
			{8'd130, 8'd45}: color_data = 12'h4a3;
			{8'd130, 8'd46}: color_data = 12'h4a3;
			{8'd130, 8'd47}: color_data = 12'h4a3;
			{8'd130, 8'd48}: color_data = 12'h4a3;
			{8'd130, 8'd49}: color_data = 12'h4a3;
			{8'd130, 8'd50}: color_data = 12'h4a3;
			{8'd130, 8'd51}: color_data = 12'h4a3;
			{8'd130, 8'd52}: color_data = 12'h4a3;
			{8'd130, 8'd53}: color_data = 12'h4a3;
			{8'd130, 8'd54}: color_data = 12'h4a3;
			{8'd130, 8'd55}: color_data = 12'h4a3;
			{8'd130, 8'd56}: color_data = 12'h4a3;
			{8'd130, 8'd57}: color_data = 12'h4a3;
			{8'd130, 8'd58}: color_data = 12'h4a3;
			{8'd130, 8'd59}: color_data = 12'h4a3;
			{8'd130, 8'd60}: color_data = 12'h4a3;
			{8'd130, 8'd61}: color_data = 12'h4a3;
			{8'd130, 8'd62}: color_data = 12'h4a3;
			{8'd130, 8'd63}: color_data = 12'h4a3;
			{8'd130, 8'd64}: color_data = 12'h4b3;
			{8'd130, 8'd65}: color_data = 12'h372;
			{8'd130, 8'd66}: color_data = 12'h000;
			{8'd130, 8'd67}: color_data = 12'h000;
			{8'd130, 8'd68}: color_data = 12'h000;
			{8'd130, 8'd69}: color_data = 12'h000;
			{8'd130, 8'd70}: color_data = 12'h000;
			{8'd130, 8'd71}: color_data = 12'h000;
			{8'd130, 8'd72}: color_data = 12'h000;
			{8'd130, 8'd100}: color_data = 12'he00;
			{8'd130, 8'd101}: color_data = 12'hf01;
			{8'd130, 8'd102}: color_data = 12'he00;
			{8'd130, 8'd103}: color_data = 12'he00;
			{8'd130, 8'd104}: color_data = 12'he00;
			{8'd130, 8'd105}: color_data = 12'he00;
			{8'd130, 8'd106}: color_data = 12'hc00;
			{8'd130, 8'd117}: color_data = 12'he00;
			{8'd130, 8'd118}: color_data = 12'he00;
			{8'd130, 8'd119}: color_data = 12'he00;
			{8'd130, 8'd120}: color_data = 12'he00;
			{8'd130, 8'd121}: color_data = 12'he00;
			{8'd130, 8'd122}: color_data = 12'he00;
			{8'd130, 8'd123}: color_data = 12'he00;
			{8'd130, 8'd127}: color_data = 12'hf00;
			{8'd130, 8'd128}: color_data = 12'he00;
			{8'd130, 8'd129}: color_data = 12'he00;
			{8'd130, 8'd130}: color_data = 12'he00;
			{8'd130, 8'd131}: color_data = 12'he00;
			{8'd130, 8'd132}: color_data = 12'he01;
			{8'd130, 8'd133}: color_data = 12'he00;
			{8'd130, 8'd138}: color_data = 12'he00;
			{8'd130, 8'd139}: color_data = 12'he00;
			{8'd130, 8'd140}: color_data = 12'he00;
			{8'd130, 8'd141}: color_data = 12'he00;
			{8'd130, 8'd142}: color_data = 12'he00;
			{8'd130, 8'd143}: color_data = 12'he01;
			{8'd130, 8'd144}: color_data = 12'he00;
			{8'd131, 8'd1}: color_data = 12'h000;
			{8'd131, 8'd2}: color_data = 12'h000;
			{8'd131, 8'd3}: color_data = 12'h540;
			{8'd131, 8'd4}: color_data = 12'hfd0;
			{8'd131, 8'd5}: color_data = 12'hfc0;
			{8'd131, 8'd6}: color_data = 12'hfc0;
			{8'd131, 8'd7}: color_data = 12'hfc0;
			{8'd131, 8'd8}: color_data = 12'hfc0;
			{8'd131, 8'd9}: color_data = 12'hfd0;
			{8'd131, 8'd10}: color_data = 12'hca0;
			{8'd131, 8'd11}: color_data = 12'h000;
			{8'd131, 8'd12}: color_data = 12'h000;
			{8'd131, 8'd13}: color_data = 12'h000;
			{8'd131, 8'd14}: color_data = 12'h000;
			{8'd131, 8'd15}: color_data = 12'h000;
			{8'd131, 8'd16}: color_data = 12'h000;
			{8'd131, 8'd17}: color_data = 12'h540;
			{8'd131, 8'd18}: color_data = 12'hfd0;
			{8'd131, 8'd19}: color_data = 12'hfc0;
			{8'd131, 8'd20}: color_data = 12'hfc0;
			{8'd131, 8'd21}: color_data = 12'hfc0;
			{8'd131, 8'd22}: color_data = 12'hfc0;
			{8'd131, 8'd23}: color_data = 12'hfd0;
			{8'd131, 8'd24}: color_data = 12'hfd0;
			{8'd131, 8'd25}: color_data = 12'h970;
			{8'd131, 8'd26}: color_data = 12'h110;
			{8'd131, 8'd27}: color_data = 12'h000;
			{8'd131, 8'd28}: color_data = 12'h000;
			{8'd131, 8'd29}: color_data = 12'h000;
			{8'd131, 8'd30}: color_data = 12'h000;
			{8'd131, 8'd31}: color_data = 12'h000;
			{8'd131, 8'd32}: color_data = 12'h000;
			{8'd131, 8'd33}: color_data = 12'h000;
			{8'd131, 8'd34}: color_data = 12'h000;
			{8'd131, 8'd35}: color_data = 12'h000;
			{8'd131, 8'd36}: color_data = 12'h000;
			{8'd131, 8'd37}: color_data = 12'h000;
			{8'd131, 8'd38}: color_data = 12'h000;
			{8'd131, 8'd39}: color_data = 12'h272;
			{8'd131, 8'd40}: color_data = 12'h4b3;
			{8'd131, 8'd41}: color_data = 12'h4b3;
			{8'd131, 8'd42}: color_data = 12'h4a3;
			{8'd131, 8'd43}: color_data = 12'h4a3;
			{8'd131, 8'd44}: color_data = 12'h4a3;
			{8'd131, 8'd45}: color_data = 12'h4a3;
			{8'd131, 8'd46}: color_data = 12'h4a3;
			{8'd131, 8'd47}: color_data = 12'h4a3;
			{8'd131, 8'd48}: color_data = 12'h4a3;
			{8'd131, 8'd49}: color_data = 12'h4a3;
			{8'd131, 8'd50}: color_data = 12'h4a3;
			{8'd131, 8'd51}: color_data = 12'h4a3;
			{8'd131, 8'd52}: color_data = 12'h4a3;
			{8'd131, 8'd53}: color_data = 12'h4a3;
			{8'd131, 8'd54}: color_data = 12'h4a3;
			{8'd131, 8'd55}: color_data = 12'h4a3;
			{8'd131, 8'd56}: color_data = 12'h4a3;
			{8'd131, 8'd57}: color_data = 12'h4a3;
			{8'd131, 8'd58}: color_data = 12'h4a3;
			{8'd131, 8'd59}: color_data = 12'h4a3;
			{8'd131, 8'd60}: color_data = 12'h4a3;
			{8'd131, 8'd61}: color_data = 12'h4a3;
			{8'd131, 8'd62}: color_data = 12'h4a3;
			{8'd131, 8'd63}: color_data = 12'h4a3;
			{8'd131, 8'd64}: color_data = 12'h4b3;
			{8'd131, 8'd65}: color_data = 12'h3a3;
			{8'd131, 8'd66}: color_data = 12'h010;
			{8'd131, 8'd67}: color_data = 12'h000;
			{8'd131, 8'd68}: color_data = 12'h000;
			{8'd131, 8'd69}: color_data = 12'h000;
			{8'd131, 8'd70}: color_data = 12'h000;
			{8'd131, 8'd71}: color_data = 12'h000;
			{8'd131, 8'd72}: color_data = 12'h000;
			{8'd131, 8'd73}: color_data = 12'h000;
			{8'd131, 8'd100}: color_data = 12'he00;
			{8'd131, 8'd101}: color_data = 12'hf01;
			{8'd131, 8'd102}: color_data = 12'he00;
			{8'd131, 8'd103}: color_data = 12'he00;
			{8'd131, 8'd104}: color_data = 12'he00;
			{8'd131, 8'd105}: color_data = 12'he00;
			{8'd131, 8'd106}: color_data = 12'hc00;
			{8'd131, 8'd117}: color_data = 12'he00;
			{8'd131, 8'd118}: color_data = 12'he01;
			{8'd131, 8'd119}: color_data = 12'he00;
			{8'd131, 8'd120}: color_data = 12'he00;
			{8'd131, 8'd121}: color_data = 12'he00;
			{8'd131, 8'd122}: color_data = 12'he01;
			{8'd131, 8'd129}: color_data = 12'he00;
			{8'd131, 8'd130}: color_data = 12'he00;
			{8'd131, 8'd131}: color_data = 12'he00;
			{8'd131, 8'd132}: color_data = 12'he00;
			{8'd131, 8'd133}: color_data = 12'he00;
			{8'd131, 8'd134}: color_data = 12'hf00;
			{8'd131, 8'd138}: color_data = 12'he00;
			{8'd131, 8'd139}: color_data = 12'he00;
			{8'd131, 8'd140}: color_data = 12'he00;
			{8'd131, 8'd141}: color_data = 12'he00;
			{8'd131, 8'd142}: color_data = 12'he00;
			{8'd131, 8'd143}: color_data = 12'he01;
			{8'd131, 8'd144}: color_data = 12'he00;
			{8'd132, 8'd1}: color_data = 12'h000;
			{8'd132, 8'd2}: color_data = 12'h000;
			{8'd132, 8'd3}: color_data = 12'h760;
			{8'd132, 8'd4}: color_data = 12'hfd0;
			{8'd132, 8'd5}: color_data = 12'hfc0;
			{8'd132, 8'd6}: color_data = 12'hfc0;
			{8'd132, 8'd7}: color_data = 12'hfc0;
			{8'd132, 8'd8}: color_data = 12'hfc0;
			{8'd132, 8'd9}: color_data = 12'hfd0;
			{8'd132, 8'd10}: color_data = 12'hfd0;
			{8'd132, 8'd11}: color_data = 12'h330;
			{8'd132, 8'd12}: color_data = 12'h000;
			{8'd132, 8'd13}: color_data = 12'h000;
			{8'd132, 8'd14}: color_data = 12'h000;
			{8'd132, 8'd15}: color_data = 12'h000;
			{8'd132, 8'd16}: color_data = 12'h000;
			{8'd132, 8'd17}: color_data = 12'h760;
			{8'd132, 8'd18}: color_data = 12'hfd0;
			{8'd132, 8'd19}: color_data = 12'hfc0;
			{8'd132, 8'd20}: color_data = 12'hfc0;
			{8'd132, 8'd21}: color_data = 12'hfc0;
			{8'd132, 8'd22}: color_data = 12'hfc0;
			{8'd132, 8'd23}: color_data = 12'hfc0;
			{8'd132, 8'd24}: color_data = 12'hfd0;
			{8'd132, 8'd25}: color_data = 12'hfd0;
			{8'd132, 8'd26}: color_data = 12'hdb0;
			{8'd132, 8'd27}: color_data = 12'h540;
			{8'd132, 8'd28}: color_data = 12'h000;
			{8'd132, 8'd29}: color_data = 12'h000;
			{8'd132, 8'd30}: color_data = 12'h000;
			{8'd132, 8'd31}: color_data = 12'h000;
			{8'd132, 8'd32}: color_data = 12'h000;
			{8'd132, 8'd33}: color_data = 12'h000;
			{8'd132, 8'd34}: color_data = 12'h000;
			{8'd132, 8'd35}: color_data = 12'h000;
			{8'd132, 8'd36}: color_data = 12'h000;
			{8'd132, 8'd37}: color_data = 12'h010;
			{8'd132, 8'd38}: color_data = 12'h382;
			{8'd132, 8'd39}: color_data = 12'h4b3;
			{8'd132, 8'd40}: color_data = 12'h4a3;
			{8'd132, 8'd41}: color_data = 12'h4a3;
			{8'd132, 8'd42}: color_data = 12'h4a3;
			{8'd132, 8'd43}: color_data = 12'h4a3;
			{8'd132, 8'd44}: color_data = 12'h4a3;
			{8'd132, 8'd45}: color_data = 12'h4a3;
			{8'd132, 8'd46}: color_data = 12'h4a3;
			{8'd132, 8'd47}: color_data = 12'h4a3;
			{8'd132, 8'd48}: color_data = 12'h4a3;
			{8'd132, 8'd49}: color_data = 12'h4a3;
			{8'd132, 8'd50}: color_data = 12'h4a3;
			{8'd132, 8'd51}: color_data = 12'h4a3;
			{8'd132, 8'd52}: color_data = 12'h4a3;
			{8'd132, 8'd53}: color_data = 12'h4a3;
			{8'd132, 8'd54}: color_data = 12'h4a3;
			{8'd132, 8'd55}: color_data = 12'h4a3;
			{8'd132, 8'd56}: color_data = 12'h4a3;
			{8'd132, 8'd57}: color_data = 12'h4a3;
			{8'd132, 8'd58}: color_data = 12'h4a3;
			{8'd132, 8'd59}: color_data = 12'h4a3;
			{8'd132, 8'd60}: color_data = 12'h4a3;
			{8'd132, 8'd61}: color_data = 12'h4a3;
			{8'd132, 8'd62}: color_data = 12'h4a3;
			{8'd132, 8'd63}: color_data = 12'h4a3;
			{8'd132, 8'd64}: color_data = 12'h4a3;
			{8'd132, 8'd65}: color_data = 12'h4b3;
			{8'd132, 8'd66}: color_data = 12'h141;
			{8'd132, 8'd67}: color_data = 12'h000;
			{8'd132, 8'd68}: color_data = 12'h000;
			{8'd132, 8'd69}: color_data = 12'h000;
			{8'd132, 8'd70}: color_data = 12'h000;
			{8'd132, 8'd71}: color_data = 12'h000;
			{8'd132, 8'd72}: color_data = 12'h000;
			{8'd132, 8'd73}: color_data = 12'h000;
			{8'd132, 8'd100}: color_data = 12'he00;
			{8'd132, 8'd101}: color_data = 12'hf01;
			{8'd132, 8'd102}: color_data = 12'he00;
			{8'd132, 8'd103}: color_data = 12'he00;
			{8'd132, 8'd104}: color_data = 12'he00;
			{8'd132, 8'd105}: color_data = 12'he00;
			{8'd132, 8'd106}: color_data = 12'hc00;
			{8'd132, 8'd117}: color_data = 12'he00;
			{8'd132, 8'd118}: color_data = 12'he01;
			{8'd132, 8'd119}: color_data = 12'he00;
			{8'd132, 8'd120}: color_data = 12'he01;
			{8'd132, 8'd121}: color_data = 12'he00;
			{8'd132, 8'd129}: color_data = 12'he00;
			{8'd132, 8'd130}: color_data = 12'he00;
			{8'd132, 8'd131}: color_data = 12'he00;
			{8'd132, 8'd132}: color_data = 12'he00;
			{8'd132, 8'd133}: color_data = 12'he00;
			{8'd132, 8'd134}: color_data = 12'hd00;
			{8'd132, 8'd138}: color_data = 12'he00;
			{8'd132, 8'd139}: color_data = 12'he00;
			{8'd132, 8'd140}: color_data = 12'he00;
			{8'd132, 8'd141}: color_data = 12'he00;
			{8'd132, 8'd142}: color_data = 12'he00;
			{8'd132, 8'd143}: color_data = 12'he01;
			{8'd132, 8'd144}: color_data = 12'he00;
			{8'd133, 8'd1}: color_data = 12'h000;
			{8'd133, 8'd2}: color_data = 12'h000;
			{8'd133, 8'd3}: color_data = 12'h320;
			{8'd133, 8'd4}: color_data = 12'hfc0;
			{8'd133, 8'd5}: color_data = 12'hfd0;
			{8'd133, 8'd6}: color_data = 12'hfc0;
			{8'd133, 8'd7}: color_data = 12'hfc0;
			{8'd133, 8'd8}: color_data = 12'hfc0;
			{8'd133, 8'd9}: color_data = 12'hfc0;
			{8'd133, 8'd10}: color_data = 12'hfd0;
			{8'd133, 8'd11}: color_data = 12'h870;
			{8'd133, 8'd12}: color_data = 12'h000;
			{8'd133, 8'd13}: color_data = 12'h110;
			{8'd133, 8'd14}: color_data = 12'h220;
			{8'd133, 8'd15}: color_data = 12'h430;
			{8'd133, 8'd16}: color_data = 12'h650;
			{8'd133, 8'd17}: color_data = 12'hca0;
			{8'd133, 8'd18}: color_data = 12'hfd0;
			{8'd133, 8'd19}: color_data = 12'hfc0;
			{8'd133, 8'd20}: color_data = 12'hfc0;
			{8'd133, 8'd21}: color_data = 12'hfc0;
			{8'd133, 8'd22}: color_data = 12'hfc0;
			{8'd133, 8'd23}: color_data = 12'hfc0;
			{8'd133, 8'd24}: color_data = 12'hfc0;
			{8'd133, 8'd25}: color_data = 12'hfc0;
			{8'd133, 8'd26}: color_data = 12'hfd0;
			{8'd133, 8'd27}: color_data = 12'hfd0;
			{8'd133, 8'd28}: color_data = 12'ha80;
			{8'd133, 8'd29}: color_data = 12'h110;
			{8'd133, 8'd30}: color_data = 12'h000;
			{8'd133, 8'd31}: color_data = 12'h000;
			{8'd133, 8'd32}: color_data = 12'h000;
			{8'd133, 8'd33}: color_data = 12'h000;
			{8'd133, 8'd34}: color_data = 12'h000;
			{8'd133, 8'd35}: color_data = 12'h000;
			{8'd133, 8'd36}: color_data = 12'h131;
			{8'd133, 8'd37}: color_data = 12'h3a3;
			{8'd133, 8'd38}: color_data = 12'h4b3;
			{8'd133, 8'd39}: color_data = 12'h4a3;
			{8'd133, 8'd40}: color_data = 12'h4a3;
			{8'd133, 8'd41}: color_data = 12'h4a3;
			{8'd133, 8'd42}: color_data = 12'h4a3;
			{8'd133, 8'd43}: color_data = 12'h4a3;
			{8'd133, 8'd44}: color_data = 12'h4a3;
			{8'd133, 8'd45}: color_data = 12'h4a3;
			{8'd133, 8'd46}: color_data = 12'h4a3;
			{8'd133, 8'd47}: color_data = 12'h4a3;
			{8'd133, 8'd48}: color_data = 12'h4a3;
			{8'd133, 8'd49}: color_data = 12'h4a3;
			{8'd133, 8'd50}: color_data = 12'h4a3;
			{8'd133, 8'd51}: color_data = 12'h4a3;
			{8'd133, 8'd52}: color_data = 12'h4a3;
			{8'd133, 8'd53}: color_data = 12'h4a3;
			{8'd133, 8'd54}: color_data = 12'h4a3;
			{8'd133, 8'd55}: color_data = 12'h4a3;
			{8'd133, 8'd56}: color_data = 12'h4a3;
			{8'd133, 8'd57}: color_data = 12'h4a3;
			{8'd133, 8'd58}: color_data = 12'h4a3;
			{8'd133, 8'd59}: color_data = 12'h4a3;
			{8'd133, 8'd60}: color_data = 12'h4a3;
			{8'd133, 8'd61}: color_data = 12'h4a3;
			{8'd133, 8'd62}: color_data = 12'h4a3;
			{8'd133, 8'd63}: color_data = 12'h4a3;
			{8'd133, 8'd64}: color_data = 12'h4a3;
			{8'd133, 8'd65}: color_data = 12'h4b3;
			{8'd133, 8'd66}: color_data = 12'h272;
			{8'd133, 8'd67}: color_data = 12'h000;
			{8'd133, 8'd68}: color_data = 12'h000;
			{8'd133, 8'd69}: color_data = 12'h000;
			{8'd133, 8'd70}: color_data = 12'h000;
			{8'd133, 8'd71}: color_data = 12'h000;
			{8'd133, 8'd72}: color_data = 12'h000;
			{8'd133, 8'd73}: color_data = 12'h000;
			{8'd133, 8'd100}: color_data = 12'he00;
			{8'd133, 8'd101}: color_data = 12'hf01;
			{8'd133, 8'd102}: color_data = 12'he00;
			{8'd133, 8'd103}: color_data = 12'he00;
			{8'd133, 8'd104}: color_data = 12'he00;
			{8'd133, 8'd105}: color_data = 12'he00;
			{8'd133, 8'd106}: color_data = 12'hc00;
			{8'd133, 8'd117}: color_data = 12'he00;
			{8'd133, 8'd118}: color_data = 12'he01;
			{8'd133, 8'd119}: color_data = 12'he00;
			{8'd133, 8'd120}: color_data = 12'he00;
			{8'd133, 8'd121}: color_data = 12'he00;
			{8'd133, 8'd122}: color_data = 12'hf00;
			{8'd133, 8'd129}: color_data = 12'he00;
			{8'd133, 8'd130}: color_data = 12'he00;
			{8'd133, 8'd131}: color_data = 12'he00;
			{8'd133, 8'd132}: color_data = 12'he00;
			{8'd133, 8'd133}: color_data = 12'he00;
			{8'd133, 8'd134}: color_data = 12'hf00;
			{8'd133, 8'd138}: color_data = 12'he00;
			{8'd133, 8'd139}: color_data = 12'he00;
			{8'd133, 8'd140}: color_data = 12'he00;
			{8'd133, 8'd141}: color_data = 12'he00;
			{8'd133, 8'd142}: color_data = 12'he00;
			{8'd133, 8'd143}: color_data = 12'he01;
			{8'd133, 8'd144}: color_data = 12'he00;
			{8'd134, 8'd1}: color_data = 12'h000;
			{8'd134, 8'd2}: color_data = 12'h000;
			{8'd134, 8'd3}: color_data = 12'h000;
			{8'd134, 8'd4}: color_data = 12'h970;
			{8'd134, 8'd5}: color_data = 12'hfd0;
			{8'd134, 8'd6}: color_data = 12'hfc0;
			{8'd134, 8'd7}: color_data = 12'hfc0;
			{8'd134, 8'd8}: color_data = 12'hfc0;
			{8'd134, 8'd9}: color_data = 12'hfc0;
			{8'd134, 8'd10}: color_data = 12'hfd0;
			{8'd134, 8'd11}: color_data = 12'hec0;
			{8'd134, 8'd12}: color_data = 12'hca0;
			{8'd134, 8'd13}: color_data = 12'heb0;
			{8'd134, 8'd14}: color_data = 12'hfc0;
			{8'd134, 8'd15}: color_data = 12'hfd0;
			{8'd134, 8'd16}: color_data = 12'hfd0;
			{8'd134, 8'd17}: color_data = 12'hfd0;
			{8'd134, 8'd18}: color_data = 12'hfc0;
			{8'd134, 8'd19}: color_data = 12'hfc0;
			{8'd134, 8'd20}: color_data = 12'hfc0;
			{8'd134, 8'd21}: color_data = 12'hfd0;
			{8'd134, 8'd22}: color_data = 12'hfc0;
			{8'd134, 8'd23}: color_data = 12'hfc0;
			{8'd134, 8'd24}: color_data = 12'hfc0;
			{8'd134, 8'd25}: color_data = 12'hfc0;
			{8'd134, 8'd26}: color_data = 12'hfc0;
			{8'd134, 8'd27}: color_data = 12'hfd0;
			{8'd134, 8'd28}: color_data = 12'hfd0;
			{8'd134, 8'd29}: color_data = 12'heb0;
			{8'd134, 8'd30}: color_data = 12'h540;
			{8'd134, 8'd31}: color_data = 12'h000;
			{8'd134, 8'd32}: color_data = 12'h000;
			{8'd134, 8'd33}: color_data = 12'h000;
			{8'd134, 8'd34}: color_data = 12'h000;
			{8'd134, 8'd35}: color_data = 12'h141;
			{8'd134, 8'd36}: color_data = 12'h4b3;
			{8'd134, 8'd37}: color_data = 12'h4b3;
			{8'd134, 8'd38}: color_data = 12'h4a3;
			{8'd134, 8'd39}: color_data = 12'h4a3;
			{8'd134, 8'd40}: color_data = 12'h4a3;
			{8'd134, 8'd41}: color_data = 12'h4a3;
			{8'd134, 8'd42}: color_data = 12'h4a3;
			{8'd134, 8'd43}: color_data = 12'h4a3;
			{8'd134, 8'd44}: color_data = 12'h4a3;
			{8'd134, 8'd45}: color_data = 12'h4a3;
			{8'd134, 8'd46}: color_data = 12'h4a3;
			{8'd134, 8'd47}: color_data = 12'h4a3;
			{8'd134, 8'd48}: color_data = 12'h4a3;
			{8'd134, 8'd49}: color_data = 12'h4a3;
			{8'd134, 8'd50}: color_data = 12'h4a3;
			{8'd134, 8'd51}: color_data = 12'h4a3;
			{8'd134, 8'd52}: color_data = 12'h4b3;
			{8'd134, 8'd53}: color_data = 12'h4b3;
			{8'd134, 8'd54}: color_data = 12'h4a3;
			{8'd134, 8'd55}: color_data = 12'h4a3;
			{8'd134, 8'd56}: color_data = 12'h4a3;
			{8'd134, 8'd57}: color_data = 12'h4a3;
			{8'd134, 8'd58}: color_data = 12'h4a3;
			{8'd134, 8'd59}: color_data = 12'h4a3;
			{8'd134, 8'd60}: color_data = 12'h4a3;
			{8'd134, 8'd61}: color_data = 12'h4a3;
			{8'd134, 8'd62}: color_data = 12'h4a3;
			{8'd134, 8'd63}: color_data = 12'h4a3;
			{8'd134, 8'd64}: color_data = 12'h4a3;
			{8'd134, 8'd65}: color_data = 12'h4b3;
			{8'd134, 8'd66}: color_data = 12'h3a3;
			{8'd134, 8'd67}: color_data = 12'h010;
			{8'd134, 8'd68}: color_data = 12'h000;
			{8'd134, 8'd69}: color_data = 12'h000;
			{8'd134, 8'd70}: color_data = 12'h000;
			{8'd134, 8'd71}: color_data = 12'h000;
			{8'd134, 8'd72}: color_data = 12'h000;
			{8'd134, 8'd73}: color_data = 12'h000;
			{8'd134, 8'd74}: color_data = 12'h000;
			{8'd134, 8'd100}: color_data = 12'he00;
			{8'd134, 8'd101}: color_data = 12'hf01;
			{8'd134, 8'd102}: color_data = 12'he00;
			{8'd134, 8'd103}: color_data = 12'he00;
			{8'd134, 8'd104}: color_data = 12'he00;
			{8'd134, 8'd105}: color_data = 12'he00;
			{8'd134, 8'd106}: color_data = 12'hc00;
			{8'd134, 8'd117}: color_data = 12'he01;
			{8'd134, 8'd118}: color_data = 12'he01;
			{8'd134, 8'd119}: color_data = 12'he00;
			{8'd134, 8'd120}: color_data = 12'he00;
			{8'd134, 8'd121}: color_data = 12'he00;
			{8'd134, 8'd122}: color_data = 12'he00;
			{8'd134, 8'd128}: color_data = 12'he00;
			{8'd134, 8'd129}: color_data = 12'he00;
			{8'd134, 8'd130}: color_data = 12'he00;
			{8'd134, 8'd131}: color_data = 12'he00;
			{8'd134, 8'd132}: color_data = 12'he00;
			{8'd134, 8'd133}: color_data = 12'he00;
			{8'd134, 8'd138}: color_data = 12'he00;
			{8'd134, 8'd139}: color_data = 12'he00;
			{8'd134, 8'd140}: color_data = 12'he00;
			{8'd134, 8'd141}: color_data = 12'he00;
			{8'd134, 8'd142}: color_data = 12'he00;
			{8'd134, 8'd143}: color_data = 12'he01;
			{8'd134, 8'd144}: color_data = 12'he00;
			{8'd135, 8'd2}: color_data = 12'h000;
			{8'd135, 8'd3}: color_data = 12'h000;
			{8'd135, 8'd4}: color_data = 12'h110;
			{8'd135, 8'd5}: color_data = 12'heb0;
			{8'd135, 8'd6}: color_data = 12'hfd0;
			{8'd135, 8'd7}: color_data = 12'hfc0;
			{8'd135, 8'd8}: color_data = 12'hfc0;
			{8'd135, 8'd9}: color_data = 12'hfc0;
			{8'd135, 8'd10}: color_data = 12'hfc0;
			{8'd135, 8'd11}: color_data = 12'hfd0;
			{8'd135, 8'd12}: color_data = 12'hfd0;
			{8'd135, 8'd13}: color_data = 12'hfd0;
			{8'd135, 8'd14}: color_data = 12'hfd0;
			{8'd135, 8'd15}: color_data = 12'hfc0;
			{8'd135, 8'd16}: color_data = 12'hfc0;
			{8'd135, 8'd17}: color_data = 12'hfc0;
			{8'd135, 8'd18}: color_data = 12'hfc0;
			{8'd135, 8'd19}: color_data = 12'hfc0;
			{8'd135, 8'd20}: color_data = 12'hfd0;
			{8'd135, 8'd21}: color_data = 12'hfd0;
			{8'd135, 8'd22}: color_data = 12'hfd0;
			{8'd135, 8'd23}: color_data = 12'hfc0;
			{8'd135, 8'd24}: color_data = 12'hfc0;
			{8'd135, 8'd25}: color_data = 12'hfc0;
			{8'd135, 8'd26}: color_data = 12'hfc0;
			{8'd135, 8'd27}: color_data = 12'hfc0;
			{8'd135, 8'd28}: color_data = 12'hfc0;
			{8'd135, 8'd29}: color_data = 12'hfd0;
			{8'd135, 8'd30}: color_data = 12'h980;
			{8'd135, 8'd31}: color_data = 12'h000;
			{8'd135, 8'd32}: color_data = 12'h000;
			{8'd135, 8'd33}: color_data = 12'h000;
			{8'd135, 8'd34}: color_data = 12'h000;
			{8'd135, 8'd35}: color_data = 12'h261;
			{8'd135, 8'd36}: color_data = 12'h4b3;
			{8'd135, 8'd37}: color_data = 12'h4a3;
			{8'd135, 8'd38}: color_data = 12'h4a3;
			{8'd135, 8'd39}: color_data = 12'h4a3;
			{8'd135, 8'd40}: color_data = 12'h4a3;
			{8'd135, 8'd41}: color_data = 12'h4a3;
			{8'd135, 8'd42}: color_data = 12'h4a3;
			{8'd135, 8'd43}: color_data = 12'h4a3;
			{8'd135, 8'd44}: color_data = 12'h4a3;
			{8'd135, 8'd45}: color_data = 12'h4a3;
			{8'd135, 8'd46}: color_data = 12'h4a3;
			{8'd135, 8'd47}: color_data = 12'h4a3;
			{8'd135, 8'd48}: color_data = 12'h4a3;
			{8'd135, 8'd49}: color_data = 12'h4a3;
			{8'd135, 8'd50}: color_data = 12'h4b3;
			{8'd135, 8'd51}: color_data = 12'h4b3;
			{8'd135, 8'd52}: color_data = 12'h4a3;
			{8'd135, 8'd53}: color_data = 12'h4a3;
			{8'd135, 8'd54}: color_data = 12'h4b3;
			{8'd135, 8'd55}: color_data = 12'h4a3;
			{8'd135, 8'd56}: color_data = 12'h4a3;
			{8'd135, 8'd57}: color_data = 12'h4a3;
			{8'd135, 8'd58}: color_data = 12'h4a3;
			{8'd135, 8'd59}: color_data = 12'h4a3;
			{8'd135, 8'd60}: color_data = 12'h4a3;
			{8'd135, 8'd61}: color_data = 12'h4a3;
			{8'd135, 8'd62}: color_data = 12'h4a3;
			{8'd135, 8'd63}: color_data = 12'h4a3;
			{8'd135, 8'd64}: color_data = 12'h4a3;
			{8'd135, 8'd65}: color_data = 12'h4a3;
			{8'd135, 8'd66}: color_data = 12'h4b3;
			{8'd135, 8'd67}: color_data = 12'h131;
			{8'd135, 8'd68}: color_data = 12'h000;
			{8'd135, 8'd69}: color_data = 12'h000;
			{8'd135, 8'd70}: color_data = 12'h000;
			{8'd135, 8'd71}: color_data = 12'h000;
			{8'd135, 8'd72}: color_data = 12'h000;
			{8'd135, 8'd73}: color_data = 12'h000;
			{8'd135, 8'd74}: color_data = 12'h000;
			{8'd135, 8'd100}: color_data = 12'he00;
			{8'd135, 8'd101}: color_data = 12'hf01;
			{8'd135, 8'd102}: color_data = 12'he00;
			{8'd135, 8'd103}: color_data = 12'he00;
			{8'd135, 8'd104}: color_data = 12'he00;
			{8'd135, 8'd105}: color_data = 12'he00;
			{8'd135, 8'd106}: color_data = 12'hc00;
			{8'd135, 8'd117}: color_data = 12'he00;
			{8'd135, 8'd118}: color_data = 12'he00;
			{8'd135, 8'd119}: color_data = 12'he00;
			{8'd135, 8'd120}: color_data = 12'he00;
			{8'd135, 8'd121}: color_data = 12'he00;
			{8'd135, 8'd122}: color_data = 12'he00;
			{8'd135, 8'd123}: color_data = 12'he00;
			{8'd135, 8'd124}: color_data = 12'he00;
			{8'd135, 8'd125}: color_data = 12'he00;
			{8'd135, 8'd126}: color_data = 12'he00;
			{8'd135, 8'd127}: color_data = 12'he00;
			{8'd135, 8'd128}: color_data = 12'he00;
			{8'd135, 8'd129}: color_data = 12'he00;
			{8'd135, 8'd130}: color_data = 12'he00;
			{8'd135, 8'd131}: color_data = 12'he00;
			{8'd135, 8'd132}: color_data = 12'hf01;
			{8'd135, 8'd133}: color_data = 12'he00;
			{8'd135, 8'd138}: color_data = 12'he00;
			{8'd135, 8'd139}: color_data = 12'he00;
			{8'd135, 8'd140}: color_data = 12'he00;
			{8'd135, 8'd141}: color_data = 12'he00;
			{8'd135, 8'd142}: color_data = 12'he00;
			{8'd135, 8'd143}: color_data = 12'he01;
			{8'd135, 8'd144}: color_data = 12'he00;
			{8'd136, 8'd2}: color_data = 12'h000;
			{8'd136, 8'd3}: color_data = 12'h000;
			{8'd136, 8'd4}: color_data = 12'h000;
			{8'd136, 8'd5}: color_data = 12'h650;
			{8'd136, 8'd6}: color_data = 12'hfd0;
			{8'd136, 8'd7}: color_data = 12'hfc0;
			{8'd136, 8'd8}: color_data = 12'hfc0;
			{8'd136, 8'd9}: color_data = 12'hfc0;
			{8'd136, 8'd10}: color_data = 12'hfc0;
			{8'd136, 8'd11}: color_data = 12'hfc0;
			{8'd136, 8'd12}: color_data = 12'hfc0;
			{8'd136, 8'd13}: color_data = 12'hfc0;
			{8'd136, 8'd14}: color_data = 12'hfc0;
			{8'd136, 8'd15}: color_data = 12'hfc0;
			{8'd136, 8'd16}: color_data = 12'hfc0;
			{8'd136, 8'd17}: color_data = 12'hfc0;
			{8'd136, 8'd18}: color_data = 12'hfc0;
			{8'd136, 8'd19}: color_data = 12'hfd0;
			{8'd136, 8'd20}: color_data = 12'hca0;
			{8'd136, 8'd21}: color_data = 12'h650;
			{8'd136, 8'd22}: color_data = 12'hfd0;
			{8'd136, 8'd23}: color_data = 12'hfd0;
			{8'd136, 8'd24}: color_data = 12'hfc0;
			{8'd136, 8'd25}: color_data = 12'hfc0;
			{8'd136, 8'd26}: color_data = 12'hfc0;
			{8'd136, 8'd27}: color_data = 12'hfc0;
			{8'd136, 8'd28}: color_data = 12'hfd0;
			{8'd136, 8'd29}: color_data = 12'hfc0;
			{8'd136, 8'd30}: color_data = 12'h330;
			{8'd136, 8'd31}: color_data = 12'h000;
			{8'd136, 8'd32}: color_data = 12'h000;
			{8'd136, 8'd33}: color_data = 12'h000;
			{8'd136, 8'd34}: color_data = 12'h000;
			{8'd136, 8'd35}: color_data = 12'h141;
			{8'd136, 8'd36}: color_data = 12'h4b3;
			{8'd136, 8'd37}: color_data = 12'h4a3;
			{8'd136, 8'd38}: color_data = 12'h4a3;
			{8'd136, 8'd39}: color_data = 12'h4a3;
			{8'd136, 8'd40}: color_data = 12'h4a3;
			{8'd136, 8'd41}: color_data = 12'h4a3;
			{8'd136, 8'd42}: color_data = 12'h4a3;
			{8'd136, 8'd43}: color_data = 12'h4a3;
			{8'd136, 8'd44}: color_data = 12'h4a3;
			{8'd136, 8'd45}: color_data = 12'h4a3;
			{8'd136, 8'd46}: color_data = 12'h4a3;
			{8'd136, 8'd47}: color_data = 12'h4a3;
			{8'd136, 8'd48}: color_data = 12'h4a3;
			{8'd136, 8'd49}: color_data = 12'h4b3;
			{8'd136, 8'd50}: color_data = 12'h4b3;
			{8'd136, 8'd51}: color_data = 12'h272;
			{8'd136, 8'd52}: color_data = 12'h010;
			{8'd136, 8'd53}: color_data = 12'h151;
			{8'd136, 8'd54}: color_data = 12'h4b3;
			{8'd136, 8'd55}: color_data = 12'h4b3;
			{8'd136, 8'd56}: color_data = 12'h4a3;
			{8'd136, 8'd57}: color_data = 12'h4a3;
			{8'd136, 8'd58}: color_data = 12'h4a3;
			{8'd136, 8'd59}: color_data = 12'h4a3;
			{8'd136, 8'd60}: color_data = 12'h4a3;
			{8'd136, 8'd61}: color_data = 12'h4a3;
			{8'd136, 8'd62}: color_data = 12'h4a3;
			{8'd136, 8'd63}: color_data = 12'h4a3;
			{8'd136, 8'd64}: color_data = 12'h4a3;
			{8'd136, 8'd65}: color_data = 12'h4a3;
			{8'd136, 8'd66}: color_data = 12'h4b3;
			{8'd136, 8'd67}: color_data = 12'h272;
			{8'd136, 8'd68}: color_data = 12'h000;
			{8'd136, 8'd69}: color_data = 12'h000;
			{8'd136, 8'd70}: color_data = 12'h000;
			{8'd136, 8'd71}: color_data = 12'h000;
			{8'd136, 8'd72}: color_data = 12'h000;
			{8'd136, 8'd73}: color_data = 12'h000;
			{8'd136, 8'd74}: color_data = 12'h000;
			{8'd136, 8'd100}: color_data = 12'he00;
			{8'd136, 8'd101}: color_data = 12'hf01;
			{8'd136, 8'd102}: color_data = 12'he00;
			{8'd136, 8'd103}: color_data = 12'he00;
			{8'd136, 8'd104}: color_data = 12'he00;
			{8'd136, 8'd105}: color_data = 12'he00;
			{8'd136, 8'd106}: color_data = 12'hf00;
			{8'd136, 8'd117}: color_data = 12'he01;
			{8'd136, 8'd118}: color_data = 12'he00;
			{8'd136, 8'd119}: color_data = 12'he00;
			{8'd136, 8'd120}: color_data = 12'he00;
			{8'd136, 8'd121}: color_data = 12'he00;
			{8'd136, 8'd122}: color_data = 12'he00;
			{8'd136, 8'd123}: color_data = 12'he00;
			{8'd136, 8'd124}: color_data = 12'he01;
			{8'd136, 8'd125}: color_data = 12'he01;
			{8'd136, 8'd126}: color_data = 12'he01;
			{8'd136, 8'd127}: color_data = 12'he01;
			{8'd136, 8'd128}: color_data = 12'he00;
			{8'd136, 8'd129}: color_data = 12'he00;
			{8'd136, 8'd130}: color_data = 12'he00;
			{8'd136, 8'd131}: color_data = 12'he00;
			{8'd136, 8'd132}: color_data = 12'he00;
			{8'd136, 8'd133}: color_data = 12'he01;
			{8'd136, 8'd138}: color_data = 12'he00;
			{8'd136, 8'd139}: color_data = 12'he00;
			{8'd136, 8'd140}: color_data = 12'he00;
			{8'd136, 8'd141}: color_data = 12'he00;
			{8'd136, 8'd142}: color_data = 12'he00;
			{8'd136, 8'd143}: color_data = 12'he01;
			{8'd136, 8'd144}: color_data = 12'he00;
			{8'd137, 8'd3}: color_data = 12'h000;
			{8'd137, 8'd4}: color_data = 12'h000;
			{8'd137, 8'd5}: color_data = 12'h000;
			{8'd137, 8'd6}: color_data = 12'hca0;
			{8'd137, 8'd7}: color_data = 12'hfd0;
			{8'd137, 8'd8}: color_data = 12'hfc0;
			{8'd137, 8'd9}: color_data = 12'hfc0;
			{8'd137, 8'd10}: color_data = 12'hfc0;
			{8'd137, 8'd11}: color_data = 12'hfc0;
			{8'd137, 8'd12}: color_data = 12'hfc0;
			{8'd137, 8'd13}: color_data = 12'hfc0;
			{8'd137, 8'd14}: color_data = 12'hfc0;
			{8'd137, 8'd15}: color_data = 12'hfc0;
			{8'd137, 8'd16}: color_data = 12'hfc0;
			{8'd137, 8'd17}: color_data = 12'hfc0;
			{8'd137, 8'd18}: color_data = 12'hfd0;
			{8'd137, 8'd19}: color_data = 12'hfd0;
			{8'd137, 8'd20}: color_data = 12'h430;
			{8'd137, 8'd21}: color_data = 12'h000;
			{8'd137, 8'd22}: color_data = 12'h760;
			{8'd137, 8'd23}: color_data = 12'hfd0;
			{8'd137, 8'd24}: color_data = 12'hfd0;
			{8'd137, 8'd25}: color_data = 12'hfc0;
			{8'd137, 8'd26}: color_data = 12'hfc0;
			{8'd137, 8'd27}: color_data = 12'hfc0;
			{8'd137, 8'd28}: color_data = 12'hfd0;
			{8'd137, 8'd29}: color_data = 12'hb90;
			{8'd137, 8'd30}: color_data = 12'h000;
			{8'd137, 8'd31}: color_data = 12'h000;
			{8'd137, 8'd32}: color_data = 12'h000;
			{8'd137, 8'd33}: color_data = 12'h000;
			{8'd137, 8'd34}: color_data = 12'h000;
			{8'd137, 8'd35}: color_data = 12'h131;
			{8'd137, 8'd36}: color_data = 12'h4b3;
			{8'd137, 8'd37}: color_data = 12'h4a3;
			{8'd137, 8'd38}: color_data = 12'h4a3;
			{8'd137, 8'd39}: color_data = 12'h4a3;
			{8'd137, 8'd40}: color_data = 12'h4a3;
			{8'd137, 8'd41}: color_data = 12'h4a3;
			{8'd137, 8'd42}: color_data = 12'h4a3;
			{8'd137, 8'd43}: color_data = 12'h4a3;
			{8'd137, 8'd44}: color_data = 12'h4a3;
			{8'd137, 8'd45}: color_data = 12'h4a3;
			{8'd137, 8'd46}: color_data = 12'h4a3;
			{8'd137, 8'd47}: color_data = 12'h4b3;
			{8'd137, 8'd48}: color_data = 12'h4b3;
			{8'd137, 8'd49}: color_data = 12'h382;
			{8'd137, 8'd50}: color_data = 12'h131;
			{8'd137, 8'd51}: color_data = 12'h000;
			{8'd137, 8'd52}: color_data = 12'h000;
			{8'd137, 8'd53}: color_data = 12'h000;
			{8'd137, 8'd54}: color_data = 12'h141;
			{8'd137, 8'd55}: color_data = 12'h4b3;
			{8'd137, 8'd56}: color_data = 12'h4b3;
			{8'd137, 8'd57}: color_data = 12'h4a3;
			{8'd137, 8'd58}: color_data = 12'h4a3;
			{8'd137, 8'd59}: color_data = 12'h4a3;
			{8'd137, 8'd60}: color_data = 12'h4a3;
			{8'd137, 8'd61}: color_data = 12'h4a3;
			{8'd137, 8'd62}: color_data = 12'h4a3;
			{8'd137, 8'd63}: color_data = 12'h4a3;
			{8'd137, 8'd64}: color_data = 12'h4a3;
			{8'd137, 8'd65}: color_data = 12'h4a3;
			{8'd137, 8'd66}: color_data = 12'h4b3;
			{8'd137, 8'd67}: color_data = 12'h393;
			{8'd137, 8'd68}: color_data = 12'h000;
			{8'd137, 8'd69}: color_data = 12'h000;
			{8'd137, 8'd70}: color_data = 12'h000;
			{8'd137, 8'd71}: color_data = 12'h000;
			{8'd137, 8'd72}: color_data = 12'h000;
			{8'd137, 8'd73}: color_data = 12'h000;
			{8'd137, 8'd74}: color_data = 12'h000;
			{8'd137, 8'd75}: color_data = 12'h000;
			{8'd137, 8'd100}: color_data = 12'he00;
			{8'd137, 8'd101}: color_data = 12'he01;
			{8'd137, 8'd102}: color_data = 12'he00;
			{8'd137, 8'd103}: color_data = 12'he00;
			{8'd137, 8'd104}: color_data = 12'he00;
			{8'd137, 8'd105}: color_data = 12'he00;
			{8'd137, 8'd106}: color_data = 12'he01;
			{8'd137, 8'd118}: color_data = 12'he00;
			{8'd137, 8'd119}: color_data = 12'hf01;
			{8'd137, 8'd120}: color_data = 12'he00;
			{8'd137, 8'd121}: color_data = 12'he00;
			{8'd137, 8'd122}: color_data = 12'he00;
			{8'd137, 8'd123}: color_data = 12'he00;
			{8'd137, 8'd124}: color_data = 12'he00;
			{8'd137, 8'd125}: color_data = 12'he00;
			{8'd137, 8'd126}: color_data = 12'he00;
			{8'd137, 8'd127}: color_data = 12'he00;
			{8'd137, 8'd128}: color_data = 12'he00;
			{8'd137, 8'd129}: color_data = 12'he00;
			{8'd137, 8'd130}: color_data = 12'he00;
			{8'd137, 8'd131}: color_data = 12'he00;
			{8'd137, 8'd132}: color_data = 12'he00;
			{8'd137, 8'd133}: color_data = 12'h700;
			{8'd137, 8'd138}: color_data = 12'he01;
			{8'd137, 8'd139}: color_data = 12'he00;
			{8'd137, 8'd140}: color_data = 12'he00;
			{8'd137, 8'd141}: color_data = 12'he00;
			{8'd137, 8'd142}: color_data = 12'he00;
			{8'd137, 8'd143}: color_data = 12'he01;
			{8'd137, 8'd144}: color_data = 12'he01;
			{8'd138, 8'd3}: color_data = 12'h000;
			{8'd138, 8'd4}: color_data = 12'h000;
			{8'd138, 8'd5}: color_data = 12'h000;
			{8'd138, 8'd6}: color_data = 12'h430;
			{8'd138, 8'd7}: color_data = 12'hfd0;
			{8'd138, 8'd8}: color_data = 12'hfd0;
			{8'd138, 8'd9}: color_data = 12'hfc0;
			{8'd138, 8'd10}: color_data = 12'hfc0;
			{8'd138, 8'd11}: color_data = 12'hfc0;
			{8'd138, 8'd12}: color_data = 12'hfc0;
			{8'd138, 8'd13}: color_data = 12'hfc0;
			{8'd138, 8'd14}: color_data = 12'hfc0;
			{8'd138, 8'd15}: color_data = 12'hfc0;
			{8'd138, 8'd16}: color_data = 12'hfc0;
			{8'd138, 8'd17}: color_data = 12'hfc0;
			{8'd138, 8'd18}: color_data = 12'hfd0;
			{8'd138, 8'd19}: color_data = 12'h980;
			{8'd138, 8'd20}: color_data = 12'h000;
			{8'd138, 8'd21}: color_data = 12'h000;
			{8'd138, 8'd22}: color_data = 12'h000;
			{8'd138, 8'd23}: color_data = 12'h980;
			{8'd138, 8'd24}: color_data = 12'hfd0;
			{8'd138, 8'd25}: color_data = 12'hfc0;
			{8'd138, 8'd26}: color_data = 12'hfc0;
			{8'd138, 8'd27}: color_data = 12'hfc0;
			{8'd138, 8'd28}: color_data = 12'hfd0;
			{8'd138, 8'd29}: color_data = 12'h540;
			{8'd138, 8'd30}: color_data = 12'h000;
			{8'd138, 8'd31}: color_data = 12'h000;
			{8'd138, 8'd32}: color_data = 12'h000;
			{8'd138, 8'd33}: color_data = 12'h000;
			{8'd138, 8'd34}: color_data = 12'h000;
			{8'd138, 8'd35}: color_data = 12'h020;
			{8'd138, 8'd36}: color_data = 12'h4a3;
			{8'd138, 8'd37}: color_data = 12'h4b3;
			{8'd138, 8'd38}: color_data = 12'h4a3;
			{8'd138, 8'd39}: color_data = 12'h4a3;
			{8'd138, 8'd40}: color_data = 12'h4a3;
			{8'd138, 8'd41}: color_data = 12'h4a3;
			{8'd138, 8'd42}: color_data = 12'h4a3;
			{8'd138, 8'd43}: color_data = 12'h4a3;
			{8'd138, 8'd44}: color_data = 12'h4a3;
			{8'd138, 8'd45}: color_data = 12'h4a3;
			{8'd138, 8'd46}: color_data = 12'h4b3;
			{8'd138, 8'd47}: color_data = 12'h3a3;
			{8'd138, 8'd48}: color_data = 12'h151;
			{8'd138, 8'd49}: color_data = 12'h000;
			{8'd138, 8'd50}: color_data = 12'h000;
			{8'd138, 8'd51}: color_data = 12'h000;
			{8'd138, 8'd52}: color_data = 12'h000;
			{8'd138, 8'd53}: color_data = 12'h000;
			{8'd138, 8'd54}: color_data = 12'h000;
			{8'd138, 8'd55}: color_data = 12'h141;
			{8'd138, 8'd56}: color_data = 12'h4a3;
			{8'd138, 8'd57}: color_data = 12'h4b3;
			{8'd138, 8'd58}: color_data = 12'h4a3;
			{8'd138, 8'd59}: color_data = 12'h4a3;
			{8'd138, 8'd60}: color_data = 12'h4a3;
			{8'd138, 8'd61}: color_data = 12'h4a3;
			{8'd138, 8'd62}: color_data = 12'h4a3;
			{8'd138, 8'd63}: color_data = 12'h4a3;
			{8'd138, 8'd64}: color_data = 12'h4a3;
			{8'd138, 8'd65}: color_data = 12'h4a3;
			{8'd138, 8'd66}: color_data = 12'h4a3;
			{8'd138, 8'd67}: color_data = 12'h4b3;
			{8'd138, 8'd68}: color_data = 12'h131;
			{8'd138, 8'd69}: color_data = 12'h000;
			{8'd138, 8'd70}: color_data = 12'h000;
			{8'd138, 8'd71}: color_data = 12'h000;
			{8'd138, 8'd72}: color_data = 12'h000;
			{8'd138, 8'd73}: color_data = 12'h000;
			{8'd138, 8'd74}: color_data = 12'h000;
			{8'd138, 8'd75}: color_data = 12'h000;
			{8'd138, 8'd100}: color_data = 12'he00;
			{8'd138, 8'd101}: color_data = 12'he01;
			{8'd138, 8'd102}: color_data = 12'he00;
			{8'd138, 8'd103}: color_data = 12'he00;
			{8'd138, 8'd104}: color_data = 12'he00;
			{8'd138, 8'd105}: color_data = 12'he00;
			{8'd138, 8'd106}: color_data = 12'he00;
			{8'd138, 8'd118}: color_data = 12'hd01;
			{8'd138, 8'd119}: color_data = 12'he00;
			{8'd138, 8'd120}: color_data = 12'hf01;
			{8'd138, 8'd121}: color_data = 12'he00;
			{8'd138, 8'd122}: color_data = 12'he00;
			{8'd138, 8'd123}: color_data = 12'he00;
			{8'd138, 8'd124}: color_data = 12'he00;
			{8'd138, 8'd125}: color_data = 12'he00;
			{8'd138, 8'd126}: color_data = 12'he00;
			{8'd138, 8'd127}: color_data = 12'he00;
			{8'd138, 8'd128}: color_data = 12'he00;
			{8'd138, 8'd129}: color_data = 12'he00;
			{8'd138, 8'd130}: color_data = 12'he00;
			{8'd138, 8'd131}: color_data = 12'he00;
			{8'd138, 8'd132}: color_data = 12'he00;
			{8'd138, 8'd138}: color_data = 12'he01;
			{8'd138, 8'd139}: color_data = 12'he00;
			{8'd138, 8'd140}: color_data = 12'he00;
			{8'd138, 8'd141}: color_data = 12'he00;
			{8'd138, 8'd142}: color_data = 12'he00;
			{8'd138, 8'd143}: color_data = 12'he00;
			{8'd138, 8'd144}: color_data = 12'he00;
			{8'd139, 8'd4}: color_data = 12'h000;
			{8'd139, 8'd5}: color_data = 12'h000;
			{8'd139, 8'd6}: color_data = 12'h000;
			{8'd139, 8'd7}: color_data = 12'ha80;
			{8'd139, 8'd8}: color_data = 12'hfd0;
			{8'd139, 8'd9}: color_data = 12'hfc0;
			{8'd139, 8'd10}: color_data = 12'hfc0;
			{8'd139, 8'd11}: color_data = 12'hfc0;
			{8'd139, 8'd12}: color_data = 12'hfc0;
			{8'd139, 8'd13}: color_data = 12'hfc0;
			{8'd139, 8'd14}: color_data = 12'hfd0;
			{8'd139, 8'd15}: color_data = 12'hfd0;
			{8'd139, 8'd16}: color_data = 12'hfd0;
			{8'd139, 8'd17}: color_data = 12'hfd0;
			{8'd139, 8'd18}: color_data = 12'heb0;
			{8'd139, 8'd19}: color_data = 12'h110;
			{8'd139, 8'd20}: color_data = 12'h000;
			{8'd139, 8'd21}: color_data = 12'h000;
			{8'd139, 8'd22}: color_data = 12'h000;
			{8'd139, 8'd23}: color_data = 12'h000;
			{8'd139, 8'd24}: color_data = 12'hb90;
			{8'd139, 8'd25}: color_data = 12'hfd0;
			{8'd139, 8'd26}: color_data = 12'hfc0;
			{8'd139, 8'd27}: color_data = 12'hfd0;
			{8'd139, 8'd28}: color_data = 12'hdb0;
			{8'd139, 8'd29}: color_data = 12'h100;
			{8'd139, 8'd30}: color_data = 12'h000;
			{8'd139, 8'd31}: color_data = 12'h000;
			{8'd139, 8'd32}: color_data = 12'h000;
			{8'd139, 8'd33}: color_data = 12'h000;
			{8'd139, 8'd34}: color_data = 12'h000;
			{8'd139, 8'd35}: color_data = 12'h010;
			{8'd139, 8'd36}: color_data = 12'h4a3;
			{8'd139, 8'd37}: color_data = 12'h4b3;
			{8'd139, 8'd38}: color_data = 12'h4a3;
			{8'd139, 8'd39}: color_data = 12'h4a3;
			{8'd139, 8'd40}: color_data = 12'h4a3;
			{8'd139, 8'd41}: color_data = 12'h4a3;
			{8'd139, 8'd42}: color_data = 12'h4a3;
			{8'd139, 8'd43}: color_data = 12'h4a3;
			{8'd139, 8'd44}: color_data = 12'h4a3;
			{8'd139, 8'd45}: color_data = 12'h4b3;
			{8'd139, 8'd46}: color_data = 12'h372;
			{8'd139, 8'd47}: color_data = 12'h010;
			{8'd139, 8'd48}: color_data = 12'h000;
			{8'd139, 8'd49}: color_data = 12'h000;
			{8'd139, 8'd50}: color_data = 12'h000;
			{8'd139, 8'd51}: color_data = 12'h000;
			{8'd139, 8'd52}: color_data = 12'h000;
			{8'd139, 8'd53}: color_data = 12'h000;
			{8'd139, 8'd54}: color_data = 12'h000;
			{8'd139, 8'd55}: color_data = 12'h000;
			{8'd139, 8'd56}: color_data = 12'h131;
			{8'd139, 8'd57}: color_data = 12'h4a3;
			{8'd139, 8'd58}: color_data = 12'h4b3;
			{8'd139, 8'd59}: color_data = 12'h4a3;
			{8'd139, 8'd60}: color_data = 12'h4a3;
			{8'd139, 8'd61}: color_data = 12'h4a3;
			{8'd139, 8'd62}: color_data = 12'h4a3;
			{8'd139, 8'd63}: color_data = 12'h4a3;
			{8'd139, 8'd64}: color_data = 12'h4a3;
			{8'd139, 8'd65}: color_data = 12'h4a3;
			{8'd139, 8'd66}: color_data = 12'h4a3;
			{8'd139, 8'd67}: color_data = 12'h4b3;
			{8'd139, 8'd68}: color_data = 12'h262;
			{8'd139, 8'd69}: color_data = 12'h000;
			{8'd139, 8'd70}: color_data = 12'h000;
			{8'd139, 8'd71}: color_data = 12'h000;
			{8'd139, 8'd72}: color_data = 12'h000;
			{8'd139, 8'd73}: color_data = 12'h000;
			{8'd139, 8'd74}: color_data = 12'h000;
			{8'd139, 8'd75}: color_data = 12'h000;
			{8'd139, 8'd100}: color_data = 12'he00;
			{8'd139, 8'd101}: color_data = 12'he01;
			{8'd139, 8'd102}: color_data = 12'he00;
			{8'd139, 8'd103}: color_data = 12'he00;
			{8'd139, 8'd104}: color_data = 12'he00;
			{8'd139, 8'd105}: color_data = 12'he00;
			{8'd139, 8'd106}: color_data = 12'he00;
			{8'd139, 8'd119}: color_data = 12'he00;
			{8'd139, 8'd120}: color_data = 12'he00;
			{8'd139, 8'd121}: color_data = 12'hf01;
			{8'd139, 8'd122}: color_data = 12'he00;
			{8'd139, 8'd123}: color_data = 12'he00;
			{8'd139, 8'd124}: color_data = 12'he00;
			{8'd139, 8'd125}: color_data = 12'he00;
			{8'd139, 8'd126}: color_data = 12'he00;
			{8'd139, 8'd127}: color_data = 12'he00;
			{8'd139, 8'd128}: color_data = 12'he00;
			{8'd139, 8'd129}: color_data = 12'he01;
			{8'd139, 8'd130}: color_data = 12'he00;
			{8'd139, 8'd131}: color_data = 12'he00;
			{8'd139, 8'd138}: color_data = 12'he00;
			{8'd139, 8'd139}: color_data = 12'he00;
			{8'd139, 8'd140}: color_data = 12'he00;
			{8'd139, 8'd141}: color_data = 12'he00;
			{8'd139, 8'd142}: color_data = 12'he00;
			{8'd139, 8'd143}: color_data = 12'he00;
			{8'd139, 8'd144}: color_data = 12'he01;
			{8'd140, 8'd5}: color_data = 12'h000;
			{8'd140, 8'd6}: color_data = 12'h000;
			{8'd140, 8'd7}: color_data = 12'h210;
			{8'd140, 8'd8}: color_data = 12'hec0;
			{8'd140, 8'd9}: color_data = 12'hfd0;
			{8'd140, 8'd10}: color_data = 12'hfd0;
			{8'd140, 8'd11}: color_data = 12'hfd0;
			{8'd140, 8'd12}: color_data = 12'hfd0;
			{8'd140, 8'd13}: color_data = 12'hfd0;
			{8'd140, 8'd14}: color_data = 12'hfc0;
			{8'd140, 8'd15}: color_data = 12'hdb0;
			{8'd140, 8'd16}: color_data = 12'hb90;
			{8'd140, 8'd17}: color_data = 12'h970;
			{8'd140, 8'd18}: color_data = 12'h330;
			{8'd140, 8'd19}: color_data = 12'h000;
			{8'd140, 8'd20}: color_data = 12'h000;
			{8'd140, 8'd21}: color_data = 12'h000;
			{8'd140, 8'd22}: color_data = 12'h000;
			{8'd140, 8'd23}: color_data = 12'h000;
			{8'd140, 8'd24}: color_data = 12'h110;
			{8'd140, 8'd25}: color_data = 12'hdb0;
			{8'd140, 8'd26}: color_data = 12'hfd0;
			{8'd140, 8'd27}: color_data = 12'hfd0;
			{8'd140, 8'd28}: color_data = 12'h860;
			{8'd140, 8'd29}: color_data = 12'h000;
			{8'd140, 8'd30}: color_data = 12'h000;
			{8'd140, 8'd31}: color_data = 12'h000;
			{8'd140, 8'd32}: color_data = 12'h000;
			{8'd140, 8'd33}: color_data = 12'h000;
			{8'd140, 8'd34}: color_data = 12'h000;
			{8'd140, 8'd35}: color_data = 12'h000;
			{8'd140, 8'd36}: color_data = 12'h392;
			{8'd140, 8'd37}: color_data = 12'h4b3;
			{8'd140, 8'd38}: color_data = 12'h4a3;
			{8'd140, 8'd39}: color_data = 12'h4a3;
			{8'd140, 8'd40}: color_data = 12'h4a3;
			{8'd140, 8'd41}: color_data = 12'h4a3;
			{8'd140, 8'd42}: color_data = 12'h4a3;
			{8'd140, 8'd43}: color_data = 12'h4a3;
			{8'd140, 8'd44}: color_data = 12'h4a3;
			{8'd140, 8'd45}: color_data = 12'h4b3;
			{8'd140, 8'd46}: color_data = 12'h262;
			{8'd140, 8'd47}: color_data = 12'h000;
			{8'd140, 8'd48}: color_data = 12'h000;
			{8'd140, 8'd49}: color_data = 12'h000;
			{8'd140, 8'd50}: color_data = 12'h000;
			{8'd140, 8'd51}: color_data = 12'h000;
			{8'd140, 8'd52}: color_data = 12'h000;
			{8'd140, 8'd53}: color_data = 12'h000;
			{8'd140, 8'd54}: color_data = 12'h000;
			{8'd140, 8'd55}: color_data = 12'h000;
			{8'd140, 8'd56}: color_data = 12'h000;
			{8'd140, 8'd57}: color_data = 12'h131;
			{8'd140, 8'd58}: color_data = 12'h3a3;
			{8'd140, 8'd59}: color_data = 12'h4b3;
			{8'd140, 8'd60}: color_data = 12'h4a3;
			{8'd140, 8'd61}: color_data = 12'h4a3;
			{8'd140, 8'd62}: color_data = 12'h4a3;
			{8'd140, 8'd63}: color_data = 12'h4a3;
			{8'd140, 8'd64}: color_data = 12'h4a3;
			{8'd140, 8'd65}: color_data = 12'h4a3;
			{8'd140, 8'd66}: color_data = 12'h4a3;
			{8'd140, 8'd67}: color_data = 12'h4b3;
			{8'd140, 8'd68}: color_data = 12'h393;
			{8'd140, 8'd69}: color_data = 12'h000;
			{8'd140, 8'd70}: color_data = 12'h000;
			{8'd140, 8'd71}: color_data = 12'h000;
			{8'd140, 8'd72}: color_data = 12'h000;
			{8'd140, 8'd73}: color_data = 12'h000;
			{8'd140, 8'd74}: color_data = 12'h000;
			{8'd140, 8'd75}: color_data = 12'h000;
			{8'd140, 8'd76}: color_data = 12'h000;
			{8'd140, 8'd100}: color_data = 12'he01;
			{8'd140, 8'd101}: color_data = 12'he00;
			{8'd140, 8'd102}: color_data = 12'he00;
			{8'd140, 8'd103}: color_data = 12'he00;
			{8'd140, 8'd104}: color_data = 12'he00;
			{8'd140, 8'd105}: color_data = 12'he00;
			{8'd140, 8'd106}: color_data = 12'he00;
			{8'd140, 8'd120}: color_data = 12'he00;
			{8'd140, 8'd121}: color_data = 12'he00;
			{8'd140, 8'd122}: color_data = 12'he00;
			{8'd140, 8'd123}: color_data = 12'he00;
			{8'd140, 8'd124}: color_data = 12'hf01;
			{8'd140, 8'd125}: color_data = 12'he01;
			{8'd140, 8'd126}: color_data = 12'he01;
			{8'd140, 8'd127}: color_data = 12'he01;
			{8'd140, 8'd128}: color_data = 12'he00;
			{8'd140, 8'd129}: color_data = 12'he00;
			{8'd140, 8'd130}: color_data = 12'he00;
			{8'd140, 8'd138}: color_data = 12'he00;
			{8'd140, 8'd139}: color_data = 12'he01;
			{8'd140, 8'd140}: color_data = 12'he00;
			{8'd140, 8'd141}: color_data = 12'he00;
			{8'd140, 8'd142}: color_data = 12'he00;
			{8'd140, 8'd143}: color_data = 12'he00;
			{8'd140, 8'd144}: color_data = 12'he00;
			{8'd141, 8'd5}: color_data = 12'h000;
			{8'd141, 8'd6}: color_data = 12'h000;
			{8'd141, 8'd7}: color_data = 12'h000;
			{8'd141, 8'd8}: color_data = 12'h750;
			{8'd141, 8'd9}: color_data = 12'hdb0;
			{8'd141, 8'd10}: color_data = 12'hb90;
			{8'd141, 8'd11}: color_data = 12'h870;
			{8'd141, 8'd12}: color_data = 12'h650;
			{8'd141, 8'd13}: color_data = 12'h430;
			{8'd141, 8'd14}: color_data = 12'h210;
			{8'd141, 8'd15}: color_data = 12'h000;
			{8'd141, 8'd16}: color_data = 12'h000;
			{8'd141, 8'd17}: color_data = 12'h000;
			{8'd141, 8'd18}: color_data = 12'h000;
			{8'd141, 8'd19}: color_data = 12'h000;
			{8'd141, 8'd20}: color_data = 12'h000;
			{8'd141, 8'd21}: color_data = 12'h000;
			{8'd141, 8'd22}: color_data = 12'h000;
			{8'd141, 8'd23}: color_data = 12'h000;
			{8'd141, 8'd24}: color_data = 12'h000;
			{8'd141, 8'd25}: color_data = 12'h320;
			{8'd141, 8'd26}: color_data = 12'hec0;
			{8'd141, 8'd27}: color_data = 12'hfc0;
			{8'd141, 8'd28}: color_data = 12'h220;
			{8'd141, 8'd29}: color_data = 12'h000;
			{8'd141, 8'd30}: color_data = 12'h000;
			{8'd141, 8'd31}: color_data = 12'h000;
			{8'd141, 8'd32}: color_data = 12'h000;
			{8'd141, 8'd33}: color_data = 12'h000;
			{8'd141, 8'd34}: color_data = 12'h000;
			{8'd141, 8'd35}: color_data = 12'h000;
			{8'd141, 8'd36}: color_data = 12'h382;
			{8'd141, 8'd37}: color_data = 12'h4b3;
			{8'd141, 8'd38}: color_data = 12'h4a3;
			{8'd141, 8'd39}: color_data = 12'h4a3;
			{8'd141, 8'd40}: color_data = 12'h4a3;
			{8'd141, 8'd41}: color_data = 12'h4a3;
			{8'd141, 8'd42}: color_data = 12'h4a3;
			{8'd141, 8'd43}: color_data = 12'h4a3;
			{8'd141, 8'd44}: color_data = 12'h4a3;
			{8'd141, 8'd45}: color_data = 12'h4b3;
			{8'd141, 8'd46}: color_data = 12'h392;
			{8'd141, 8'd47}: color_data = 12'h000;
			{8'd141, 8'd48}: color_data = 12'h000;
			{8'd141, 8'd49}: color_data = 12'h000;
			{8'd141, 8'd50}: color_data = 12'h000;
			{8'd141, 8'd51}: color_data = 12'h000;
			{8'd141, 8'd52}: color_data = 12'h000;
			{8'd141, 8'd53}: color_data = 12'h000;
			{8'd141, 8'd54}: color_data = 12'h000;
			{8'd141, 8'd55}: color_data = 12'h000;
			{8'd141, 8'd56}: color_data = 12'h000;
			{8'd141, 8'd57}: color_data = 12'h000;
			{8'd141, 8'd58}: color_data = 12'h382;
			{8'd141, 8'd59}: color_data = 12'h4b3;
			{8'd141, 8'd60}: color_data = 12'h4a3;
			{8'd141, 8'd61}: color_data = 12'h4a3;
			{8'd141, 8'd62}: color_data = 12'h4a3;
			{8'd141, 8'd63}: color_data = 12'h4a3;
			{8'd141, 8'd64}: color_data = 12'h4a3;
			{8'd141, 8'd65}: color_data = 12'h4a3;
			{8'd141, 8'd66}: color_data = 12'h4a3;
			{8'd141, 8'd67}: color_data = 12'h4a3;
			{8'd141, 8'd68}: color_data = 12'h4b3;
			{8'd141, 8'd69}: color_data = 12'h131;
			{8'd141, 8'd70}: color_data = 12'h000;
			{8'd141, 8'd71}: color_data = 12'h000;
			{8'd141, 8'd72}: color_data = 12'h000;
			{8'd141, 8'd73}: color_data = 12'h000;
			{8'd141, 8'd74}: color_data = 12'h000;
			{8'd141, 8'd75}: color_data = 12'h000;
			{8'd141, 8'd76}: color_data = 12'h000;
			{8'd141, 8'd100}: color_data = 12'he01;
			{8'd141, 8'd101}: color_data = 12'he00;
			{8'd141, 8'd102}: color_data = 12'he00;
			{8'd141, 8'd103}: color_data = 12'he00;
			{8'd141, 8'd104}: color_data = 12'he00;
			{8'd141, 8'd105}: color_data = 12'he01;
			{8'd141, 8'd106}: color_data = 12'he00;
			{8'd141, 8'd122}: color_data = 12'he00;
			{8'd141, 8'd123}: color_data = 12'he01;
			{8'd141, 8'd124}: color_data = 12'he00;
			{8'd141, 8'd125}: color_data = 12'he00;
			{8'd141, 8'd126}: color_data = 12'he00;
			{8'd141, 8'd127}: color_data = 12'he00;
			{8'd141, 8'd128}: color_data = 12'he00;
			{8'd141, 8'd129}: color_data = 12'hf00;
			{8'd141, 8'd138}: color_data = 12'he00;
			{8'd141, 8'd139}: color_data = 12'he00;
			{8'd141, 8'd140}: color_data = 12'he00;
			{8'd141, 8'd141}: color_data = 12'he00;
			{8'd141, 8'd142}: color_data = 12'he00;
			{8'd141, 8'd143}: color_data = 12'he00;
			{8'd141, 8'd144}: color_data = 12'hf00;
			{8'd142, 8'd6}: color_data = 12'h000;
			{8'd142, 8'd7}: color_data = 12'h000;
			{8'd142, 8'd8}: color_data = 12'h000;
			{8'd142, 8'd9}: color_data = 12'h000;
			{8'd142, 8'd10}: color_data = 12'h000;
			{8'd142, 8'd11}: color_data = 12'h000;
			{8'd142, 8'd12}: color_data = 12'h000;
			{8'd142, 8'd13}: color_data = 12'h000;
			{8'd142, 8'd14}: color_data = 12'h000;
			{8'd142, 8'd15}: color_data = 12'h000;
			{8'd142, 8'd16}: color_data = 12'h000;
			{8'd142, 8'd17}: color_data = 12'h000;
			{8'd142, 8'd18}: color_data = 12'h000;
			{8'd142, 8'd19}: color_data = 12'h000;
			{8'd142, 8'd20}: color_data = 12'h000;
			{8'd142, 8'd21}: color_data = 12'h000;
			{8'd142, 8'd22}: color_data = 12'h000;
			{8'd142, 8'd23}: color_data = 12'h000;
			{8'd142, 8'd24}: color_data = 12'h000;
			{8'd142, 8'd25}: color_data = 12'h000;
			{8'd142, 8'd26}: color_data = 12'h540;
			{8'd142, 8'd27}: color_data = 12'h970;
			{8'd142, 8'd28}: color_data = 12'h000;
			{8'd142, 8'd29}: color_data = 12'h000;
			{8'd142, 8'd30}: color_data = 12'h000;
			{8'd142, 8'd31}: color_data = 12'h000;
			{8'd142, 8'd32}: color_data = 12'h000;
			{8'd142, 8'd33}: color_data = 12'h000;
			{8'd142, 8'd34}: color_data = 12'h000;
			{8'd142, 8'd35}: color_data = 12'h000;
			{8'd142, 8'd36}: color_data = 12'h372;
			{8'd142, 8'd37}: color_data = 12'h4b3;
			{8'd142, 8'd38}: color_data = 12'h4a3;
			{8'd142, 8'd39}: color_data = 12'h4a3;
			{8'd142, 8'd40}: color_data = 12'h4a3;
			{8'd142, 8'd41}: color_data = 12'h4a3;
			{8'd142, 8'd42}: color_data = 12'h4a3;
			{8'd142, 8'd43}: color_data = 12'h4a3;
			{8'd142, 8'd44}: color_data = 12'h4a3;
			{8'd142, 8'd45}: color_data = 12'h4b3;
			{8'd142, 8'd46}: color_data = 12'h4a3;
			{8'd142, 8'd47}: color_data = 12'h020;
			{8'd142, 8'd48}: color_data = 12'h000;
			{8'd142, 8'd49}: color_data = 12'h000;
			{8'd142, 8'd50}: color_data = 12'h000;
			{8'd142, 8'd51}: color_data = 12'h000;
			{8'd142, 8'd52}: color_data = 12'h000;
			{8'd142, 8'd53}: color_data = 12'h000;
			{8'd142, 8'd54}: color_data = 12'h000;
			{8'd142, 8'd55}: color_data = 12'h000;
			{8'd142, 8'd56}: color_data = 12'h000;
			{8'd142, 8'd57}: color_data = 12'h130;
			{8'd142, 8'd58}: color_data = 12'h4a3;
			{8'd142, 8'd59}: color_data = 12'h4b3;
			{8'd142, 8'd60}: color_data = 12'h4a3;
			{8'd142, 8'd61}: color_data = 12'h4a3;
			{8'd142, 8'd62}: color_data = 12'h4a3;
			{8'd142, 8'd63}: color_data = 12'h4a3;
			{8'd142, 8'd64}: color_data = 12'h4a3;
			{8'd142, 8'd65}: color_data = 12'h4a3;
			{8'd142, 8'd66}: color_data = 12'h4a3;
			{8'd142, 8'd67}: color_data = 12'h4a3;
			{8'd142, 8'd68}: color_data = 12'h4b3;
			{8'd142, 8'd69}: color_data = 12'h261;
			{8'd142, 8'd70}: color_data = 12'h000;
			{8'd142, 8'd71}: color_data = 12'h000;
			{8'd142, 8'd72}: color_data = 12'h000;
			{8'd142, 8'd73}: color_data = 12'h000;
			{8'd142, 8'd74}: color_data = 12'h000;
			{8'd142, 8'd75}: color_data = 12'h000;
			{8'd142, 8'd76}: color_data = 12'h000;
			{8'd142, 8'd101}: color_data = 12'he00;
			{8'd142, 8'd102}: color_data = 12'he00;
			{8'd142, 8'd103}: color_data = 12'he00;
			{8'd142, 8'd104}: color_data = 12'he00;
			{8'd142, 8'd105}: color_data = 12'he00;
			{8'd142, 8'd106}: color_data = 12'he00;
			{8'd142, 8'd107}: color_data = 12'he01;
			{8'd142, 8'd137}: color_data = 12'he00;
			{8'd142, 8'd138}: color_data = 12'he00;
			{8'd142, 8'd139}: color_data = 12'he00;
			{8'd142, 8'd140}: color_data = 12'he00;
			{8'd142, 8'd141}: color_data = 12'he00;
			{8'd142, 8'd142}: color_data = 12'he01;
			{8'd142, 8'd143}: color_data = 12'he00;
			{8'd143, 8'd6}: color_data = 12'h000;
			{8'd143, 8'd7}: color_data = 12'h000;
			{8'd143, 8'd8}: color_data = 12'h000;
			{8'd143, 8'd9}: color_data = 12'h000;
			{8'd143, 8'd10}: color_data = 12'h000;
			{8'd143, 8'd11}: color_data = 12'h000;
			{8'd143, 8'd12}: color_data = 12'h000;
			{8'd143, 8'd13}: color_data = 12'h000;
			{8'd143, 8'd14}: color_data = 12'h000;
			{8'd143, 8'd15}: color_data = 12'h000;
			{8'd143, 8'd16}: color_data = 12'h000;
			{8'd143, 8'd17}: color_data = 12'h000;
			{8'd143, 8'd18}: color_data = 12'h000;
			{8'd143, 8'd19}: color_data = 12'h000;
			{8'd143, 8'd20}: color_data = 12'h000;
			{8'd143, 8'd21}: color_data = 12'h000;
			{8'd143, 8'd24}: color_data = 12'h000;
			{8'd143, 8'd25}: color_data = 12'h000;
			{8'd143, 8'd26}: color_data = 12'h000;
			{8'd143, 8'd27}: color_data = 12'h000;
			{8'd143, 8'd28}: color_data = 12'h000;
			{8'd143, 8'd29}: color_data = 12'h000;
			{8'd143, 8'd30}: color_data = 12'h000;
			{8'd143, 8'd31}: color_data = 12'h000;
			{8'd143, 8'd32}: color_data = 12'h000;
			{8'd143, 8'd33}: color_data = 12'h000;
			{8'd143, 8'd34}: color_data = 12'h000;
			{8'd143, 8'd35}: color_data = 12'h000;
			{8'd143, 8'd36}: color_data = 12'h261;
			{8'd143, 8'd37}: color_data = 12'h4b3;
			{8'd143, 8'd38}: color_data = 12'h4a3;
			{8'd143, 8'd39}: color_data = 12'h4a3;
			{8'd143, 8'd40}: color_data = 12'h4a3;
			{8'd143, 8'd41}: color_data = 12'h4a3;
			{8'd143, 8'd42}: color_data = 12'h4a3;
			{8'd143, 8'd43}: color_data = 12'h4a3;
			{8'd143, 8'd44}: color_data = 12'h4a3;
			{8'd143, 8'd45}: color_data = 12'h4a3;
			{8'd143, 8'd46}: color_data = 12'h4b3;
			{8'd143, 8'd47}: color_data = 12'h141;
			{8'd143, 8'd48}: color_data = 12'h000;
			{8'd143, 8'd49}: color_data = 12'h000;
			{8'd143, 8'd50}: color_data = 12'h000;
			{8'd143, 8'd51}: color_data = 12'h000;
			{8'd143, 8'd52}: color_data = 12'h000;
			{8'd143, 8'd53}: color_data = 12'h000;
			{8'd143, 8'd54}: color_data = 12'h000;
			{8'd143, 8'd55}: color_data = 12'h000;
			{8'd143, 8'd56}: color_data = 12'h000;
			{8'd143, 8'd57}: color_data = 12'h372;
			{8'd143, 8'd58}: color_data = 12'h4b3;
			{8'd143, 8'd59}: color_data = 12'h4a3;
			{8'd143, 8'd60}: color_data = 12'h4a3;
			{8'd143, 8'd61}: color_data = 12'h4a3;
			{8'd143, 8'd62}: color_data = 12'h4a3;
			{8'd143, 8'd63}: color_data = 12'h4a3;
			{8'd143, 8'd64}: color_data = 12'h4a3;
			{8'd143, 8'd65}: color_data = 12'h4a3;
			{8'd143, 8'd66}: color_data = 12'h4a3;
			{8'd143, 8'd67}: color_data = 12'h4a3;
			{8'd143, 8'd68}: color_data = 12'h4b3;
			{8'd143, 8'd69}: color_data = 12'h151;
			{8'd143, 8'd70}: color_data = 12'h000;
			{8'd143, 8'd71}: color_data = 12'h000;
			{8'd143, 8'd72}: color_data = 12'h000;
			{8'd143, 8'd73}: color_data = 12'h000;
			{8'd143, 8'd74}: color_data = 12'h000;
			{8'd143, 8'd75}: color_data = 12'h000;
			{8'd143, 8'd76}: color_data = 12'h000;
			{8'd143, 8'd101}: color_data = 12'he01;
			{8'd143, 8'd102}: color_data = 12'he01;
			{8'd143, 8'd103}: color_data = 12'he00;
			{8'd143, 8'd104}: color_data = 12'he00;
			{8'd143, 8'd105}: color_data = 12'he00;
			{8'd143, 8'd106}: color_data = 12'he00;
			{8'd143, 8'd107}: color_data = 12'he00;
			{8'd143, 8'd137}: color_data = 12'he00;
			{8'd143, 8'd138}: color_data = 12'he00;
			{8'd143, 8'd139}: color_data = 12'he00;
			{8'd143, 8'd140}: color_data = 12'he00;
			{8'd143, 8'd141}: color_data = 12'he00;
			{8'd143, 8'd142}: color_data = 12'he00;
			{8'd143, 8'd143}: color_data = 12'he00;
			{8'd144, 8'd7}: color_data = 12'h000;
			{8'd144, 8'd8}: color_data = 12'h000;
			{8'd144, 8'd9}: color_data = 12'h000;
			{8'd144, 8'd10}: color_data = 12'h000;
			{8'd144, 8'd11}: color_data = 12'h000;
			{8'd144, 8'd12}: color_data = 12'h000;
			{8'd144, 8'd13}: color_data = 12'h000;
			{8'd144, 8'd14}: color_data = 12'h000;
			{8'd144, 8'd15}: color_data = 12'h000;
			{8'd144, 8'd25}: color_data = 12'h000;
			{8'd144, 8'd26}: color_data = 12'h000;
			{8'd144, 8'd27}: color_data = 12'h000;
			{8'd144, 8'd28}: color_data = 12'h000;
			{8'd144, 8'd29}: color_data = 12'h000;
			{8'd144, 8'd30}: color_data = 12'h000;
			{8'd144, 8'd31}: color_data = 12'h000;
			{8'd144, 8'd32}: color_data = 12'h000;
			{8'd144, 8'd33}: color_data = 12'h000;
			{8'd144, 8'd34}: color_data = 12'h000;
			{8'd144, 8'd35}: color_data = 12'h000;
			{8'd144, 8'd36}: color_data = 12'h251;
			{8'd144, 8'd37}: color_data = 12'h4b3;
			{8'd144, 8'd38}: color_data = 12'h4a3;
			{8'd144, 8'd39}: color_data = 12'h4a3;
			{8'd144, 8'd40}: color_data = 12'h4a3;
			{8'd144, 8'd41}: color_data = 12'h4a3;
			{8'd144, 8'd42}: color_data = 12'h4a3;
			{8'd144, 8'd43}: color_data = 12'h4a3;
			{8'd144, 8'd44}: color_data = 12'h4a3;
			{8'd144, 8'd45}: color_data = 12'h4a3;
			{8'd144, 8'd46}: color_data = 12'h4b3;
			{8'd144, 8'd47}: color_data = 12'h372;
			{8'd144, 8'd48}: color_data = 12'h000;
			{8'd144, 8'd49}: color_data = 12'h000;
			{8'd144, 8'd50}: color_data = 12'h000;
			{8'd144, 8'd51}: color_data = 12'h000;
			{8'd144, 8'd52}: color_data = 12'h000;
			{8'd144, 8'd53}: color_data = 12'h000;
			{8'd144, 8'd54}: color_data = 12'h000;
			{8'd144, 8'd55}: color_data = 12'h000;
			{8'd144, 8'd56}: color_data = 12'h120;
			{8'd144, 8'd57}: color_data = 12'h4b3;
			{8'd144, 8'd58}: color_data = 12'h4b3;
			{8'd144, 8'd59}: color_data = 12'h4a3;
			{8'd144, 8'd60}: color_data = 12'h4a3;
			{8'd144, 8'd61}: color_data = 12'h4a3;
			{8'd144, 8'd62}: color_data = 12'h4a3;
			{8'd144, 8'd63}: color_data = 12'h4a3;
			{8'd144, 8'd64}: color_data = 12'h4a3;
			{8'd144, 8'd65}: color_data = 12'h4a3;
			{8'd144, 8'd66}: color_data = 12'h4a3;
			{8'd144, 8'd67}: color_data = 12'h4b3;
			{8'd144, 8'd68}: color_data = 12'h3a3;
			{8'd144, 8'd69}: color_data = 12'h010;
			{8'd144, 8'd70}: color_data = 12'h000;
			{8'd144, 8'd71}: color_data = 12'h000;
			{8'd144, 8'd72}: color_data = 12'h000;
			{8'd144, 8'd73}: color_data = 12'h000;
			{8'd144, 8'd74}: color_data = 12'h000;
			{8'd144, 8'd75}: color_data = 12'h000;
			{8'd144, 8'd76}: color_data = 12'h000;
			{8'd144, 8'd101}: color_data = 12'he01;
			{8'd144, 8'd102}: color_data = 12'he00;
			{8'd144, 8'd103}: color_data = 12'he00;
			{8'd144, 8'd104}: color_data = 12'he00;
			{8'd144, 8'd105}: color_data = 12'he00;
			{8'd144, 8'd106}: color_data = 12'he00;
			{8'd144, 8'd107}: color_data = 12'he00;
			{8'd144, 8'd108}: color_data = 12'hc00;
			{8'd144, 8'd136}: color_data = 12'he00;
			{8'd144, 8'd137}: color_data = 12'he00;
			{8'd144, 8'd138}: color_data = 12'he00;
			{8'd144, 8'd139}: color_data = 12'he00;
			{8'd144, 8'd140}: color_data = 12'he00;
			{8'd144, 8'd141}: color_data = 12'he00;
			{8'd144, 8'd142}: color_data = 12'he00;
			{8'd144, 8'd143}: color_data = 12'he00;
			{8'd145, 8'd25}: color_data = 12'h000;
			{8'd145, 8'd26}: color_data = 12'h000;
			{8'd145, 8'd27}: color_data = 12'h000;
			{8'd145, 8'd28}: color_data = 12'h000;
			{8'd145, 8'd29}: color_data = 12'h000;
			{8'd145, 8'd30}: color_data = 12'h000;
			{8'd145, 8'd31}: color_data = 12'h000;
			{8'd145, 8'd32}: color_data = 12'h000;
			{8'd145, 8'd33}: color_data = 12'h000;
			{8'd145, 8'd34}: color_data = 12'h000;
			{8'd145, 8'd35}: color_data = 12'h000;
			{8'd145, 8'd36}: color_data = 12'h131;
			{8'd145, 8'd37}: color_data = 12'h4b3;
			{8'd145, 8'd38}: color_data = 12'h4a3;
			{8'd145, 8'd39}: color_data = 12'h4a3;
			{8'd145, 8'd40}: color_data = 12'h4a3;
			{8'd145, 8'd41}: color_data = 12'h4a3;
			{8'd145, 8'd42}: color_data = 12'h4a3;
			{8'd145, 8'd43}: color_data = 12'h4a3;
			{8'd145, 8'd44}: color_data = 12'h4a3;
			{8'd145, 8'd45}: color_data = 12'h4a3;
			{8'd145, 8'd46}: color_data = 12'h4b3;
			{8'd145, 8'd47}: color_data = 12'h393;
			{8'd145, 8'd48}: color_data = 12'h000;
			{8'd145, 8'd49}: color_data = 12'h000;
			{8'd145, 8'd50}: color_data = 12'h000;
			{8'd145, 8'd51}: color_data = 12'h000;
			{8'd145, 8'd52}: color_data = 12'h000;
			{8'd145, 8'd53}: color_data = 12'h000;
			{8'd145, 8'd54}: color_data = 12'h000;
			{8'd145, 8'd55}: color_data = 12'h000;
			{8'd145, 8'd56}: color_data = 12'h372;
			{8'd145, 8'd57}: color_data = 12'h4b3;
			{8'd145, 8'd58}: color_data = 12'h4a3;
			{8'd145, 8'd59}: color_data = 12'h4a3;
			{8'd145, 8'd60}: color_data = 12'h4a3;
			{8'd145, 8'd61}: color_data = 12'h4a3;
			{8'd145, 8'd62}: color_data = 12'h4a3;
			{8'd145, 8'd63}: color_data = 12'h4a3;
			{8'd145, 8'd64}: color_data = 12'h4a3;
			{8'd145, 8'd65}: color_data = 12'h4a3;
			{8'd145, 8'd66}: color_data = 12'h4a3;
			{8'd145, 8'd67}: color_data = 12'h4b3;
			{8'd145, 8'd68}: color_data = 12'h261;
			{8'd145, 8'd69}: color_data = 12'h000;
			{8'd145, 8'd70}: color_data = 12'h000;
			{8'd145, 8'd71}: color_data = 12'h000;
			{8'd145, 8'd72}: color_data = 12'h000;
			{8'd145, 8'd73}: color_data = 12'h000;
			{8'd145, 8'd74}: color_data = 12'h000;
			{8'd145, 8'd75}: color_data = 12'h000;
			{8'd145, 8'd102}: color_data = 12'he00;
			{8'd145, 8'd103}: color_data = 12'he00;
			{8'd145, 8'd104}: color_data = 12'he00;
			{8'd145, 8'd105}: color_data = 12'he00;
			{8'd145, 8'd106}: color_data = 12'he00;
			{8'd145, 8'd107}: color_data = 12'he00;
			{8'd145, 8'd108}: color_data = 12'he00;
			{8'd145, 8'd136}: color_data = 12'he00;
			{8'd145, 8'd137}: color_data = 12'he00;
			{8'd145, 8'd138}: color_data = 12'he00;
			{8'd145, 8'd139}: color_data = 12'he00;
			{8'd145, 8'd140}: color_data = 12'he00;
			{8'd145, 8'd141}: color_data = 12'he01;
			{8'd145, 8'd142}: color_data = 12'he00;
			{8'd146, 8'd26}: color_data = 12'h000;
			{8'd146, 8'd27}: color_data = 12'h000;
			{8'd146, 8'd28}: color_data = 12'h000;
			{8'd146, 8'd29}: color_data = 12'h000;
			{8'd146, 8'd30}: color_data = 12'h000;
			{8'd146, 8'd31}: color_data = 12'h000;
			{8'd146, 8'd33}: color_data = 12'h000;
			{8'd146, 8'd34}: color_data = 12'h000;
			{8'd146, 8'd35}: color_data = 12'h000;
			{8'd146, 8'd36}: color_data = 12'h120;
			{8'd146, 8'd37}: color_data = 12'h4b3;
			{8'd146, 8'd38}: color_data = 12'h4b3;
			{8'd146, 8'd39}: color_data = 12'h4a3;
			{8'd146, 8'd40}: color_data = 12'h4a3;
			{8'd146, 8'd41}: color_data = 12'h4a3;
			{8'd146, 8'd42}: color_data = 12'h4a3;
			{8'd146, 8'd43}: color_data = 12'h4a3;
			{8'd146, 8'd44}: color_data = 12'h4a3;
			{8'd146, 8'd45}: color_data = 12'h4a3;
			{8'd146, 8'd46}: color_data = 12'h4a3;
			{8'd146, 8'd47}: color_data = 12'h4b3;
			{8'd146, 8'd48}: color_data = 12'h251;
			{8'd146, 8'd49}: color_data = 12'h020;
			{8'd146, 8'd50}: color_data = 12'h010;
			{8'd146, 8'd51}: color_data = 12'h000;
			{8'd146, 8'd52}: color_data = 12'h000;
			{8'd146, 8'd53}: color_data = 12'h000;
			{8'd146, 8'd54}: color_data = 12'h000;
			{8'd146, 8'd55}: color_data = 12'h120;
			{8'd146, 8'd56}: color_data = 12'h4b3;
			{8'd146, 8'd57}: color_data = 12'h4b3;
			{8'd146, 8'd58}: color_data = 12'h4a3;
			{8'd146, 8'd59}: color_data = 12'h4a3;
			{8'd146, 8'd60}: color_data = 12'h4a3;
			{8'd146, 8'd61}: color_data = 12'h4a3;
			{8'd146, 8'd62}: color_data = 12'h4a3;
			{8'd146, 8'd63}: color_data = 12'h4a3;
			{8'd146, 8'd64}: color_data = 12'h4a3;
			{8'd146, 8'd65}: color_data = 12'h4a3;
			{8'd146, 8'd66}: color_data = 12'h4b3;
			{8'd146, 8'd67}: color_data = 12'h4a3;
			{8'd146, 8'd68}: color_data = 12'h010;
			{8'd146, 8'd69}: color_data = 12'h000;
			{8'd146, 8'd70}: color_data = 12'h000;
			{8'd146, 8'd71}: color_data = 12'h000;
			{8'd146, 8'd72}: color_data = 12'h000;
			{8'd146, 8'd73}: color_data = 12'h000;
			{8'd146, 8'd74}: color_data = 12'h000;
			{8'd146, 8'd75}: color_data = 12'h000;
			{8'd146, 8'd102}: color_data = 12'he00;
			{8'd146, 8'd103}: color_data = 12'he00;
			{8'd146, 8'd104}: color_data = 12'he00;
			{8'd146, 8'd105}: color_data = 12'he00;
			{8'd146, 8'd106}: color_data = 12'he00;
			{8'd146, 8'd107}: color_data = 12'he00;
			{8'd146, 8'd108}: color_data = 12'he00;
			{8'd146, 8'd109}: color_data = 12'he00;
			{8'd146, 8'd135}: color_data = 12'he00;
			{8'd146, 8'd136}: color_data = 12'he00;
			{8'd146, 8'd137}: color_data = 12'he00;
			{8'd146, 8'd138}: color_data = 12'he00;
			{8'd146, 8'd139}: color_data = 12'he00;
			{8'd146, 8'd140}: color_data = 12'he00;
			{8'd146, 8'd141}: color_data = 12'he00;
			{8'd146, 8'd142}: color_data = 12'he01;
			{8'd147, 8'd34}: color_data = 12'h000;
			{8'd147, 8'd35}: color_data = 12'h000;
			{8'd147, 8'd36}: color_data = 12'h010;
			{8'd147, 8'd37}: color_data = 12'h4a3;
			{8'd147, 8'd38}: color_data = 12'h4b3;
			{8'd147, 8'd39}: color_data = 12'h4a3;
			{8'd147, 8'd40}: color_data = 12'h4a3;
			{8'd147, 8'd41}: color_data = 12'h4a3;
			{8'd147, 8'd42}: color_data = 12'h4a3;
			{8'd147, 8'd43}: color_data = 12'h4a3;
			{8'd147, 8'd44}: color_data = 12'h4a3;
			{8'd147, 8'd45}: color_data = 12'h4a3;
			{8'd147, 8'd46}: color_data = 12'h4a3;
			{8'd147, 8'd47}: color_data = 12'h4a3;
			{8'd147, 8'd48}: color_data = 12'h4b3;
			{8'd147, 8'd49}: color_data = 12'h4b3;
			{8'd147, 8'd50}: color_data = 12'h4a3;
			{8'd147, 8'd51}: color_data = 12'h393;
			{8'd147, 8'd52}: color_data = 12'h382;
			{8'd147, 8'd53}: color_data = 12'h372;
			{8'd147, 8'd54}: color_data = 12'h261;
			{8'd147, 8'd55}: color_data = 12'h382;
			{8'd147, 8'd56}: color_data = 12'h4b3;
			{8'd147, 8'd57}: color_data = 12'h4a3;
			{8'd147, 8'd58}: color_data = 12'h4a3;
			{8'd147, 8'd59}: color_data = 12'h4a3;
			{8'd147, 8'd60}: color_data = 12'h4a3;
			{8'd147, 8'd61}: color_data = 12'h4a3;
			{8'd147, 8'd62}: color_data = 12'h4a3;
			{8'd147, 8'd63}: color_data = 12'h4a3;
			{8'd147, 8'd64}: color_data = 12'h4a3;
			{8'd147, 8'd65}: color_data = 12'h4a3;
			{8'd147, 8'd66}: color_data = 12'h4b3;
			{8'd147, 8'd67}: color_data = 12'h262;
			{8'd147, 8'd68}: color_data = 12'h000;
			{8'd147, 8'd69}: color_data = 12'h000;
			{8'd147, 8'd70}: color_data = 12'h000;
			{8'd147, 8'd71}: color_data = 12'h000;
			{8'd147, 8'd72}: color_data = 12'h000;
			{8'd147, 8'd73}: color_data = 12'h000;
			{8'd147, 8'd74}: color_data = 12'h000;
			{8'd147, 8'd102}: color_data = 12'ha00;
			{8'd147, 8'd103}: color_data = 12'he00;
			{8'd147, 8'd104}: color_data = 12'he01;
			{8'd147, 8'd105}: color_data = 12'he00;
			{8'd147, 8'd106}: color_data = 12'he00;
			{8'd147, 8'd107}: color_data = 12'he00;
			{8'd147, 8'd108}: color_data = 12'he00;
			{8'd147, 8'd109}: color_data = 12'he00;
			{8'd147, 8'd110}: color_data = 12'he01;
			{8'd147, 8'd134}: color_data = 12'he00;
			{8'd147, 8'd135}: color_data = 12'he00;
			{8'd147, 8'd136}: color_data = 12'he00;
			{8'd147, 8'd137}: color_data = 12'he00;
			{8'd147, 8'd138}: color_data = 12'he00;
			{8'd147, 8'd139}: color_data = 12'he00;
			{8'd147, 8'd140}: color_data = 12'hf01;
			{8'd147, 8'd141}: color_data = 12'he00;
			{8'd148, 8'd34}: color_data = 12'h000;
			{8'd148, 8'd35}: color_data = 12'h000;
			{8'd148, 8'd36}: color_data = 12'h000;
			{8'd148, 8'd37}: color_data = 12'h393;
			{8'd148, 8'd38}: color_data = 12'h4b3;
			{8'd148, 8'd39}: color_data = 12'h4a3;
			{8'd148, 8'd40}: color_data = 12'h4a3;
			{8'd148, 8'd41}: color_data = 12'h4a3;
			{8'd148, 8'd42}: color_data = 12'h4a3;
			{8'd148, 8'd43}: color_data = 12'h4a3;
			{8'd148, 8'd44}: color_data = 12'h4a3;
			{8'd148, 8'd45}: color_data = 12'h4a3;
			{8'd148, 8'd46}: color_data = 12'h4a3;
			{8'd148, 8'd47}: color_data = 12'h4a3;
			{8'd148, 8'd48}: color_data = 12'h4a3;
			{8'd148, 8'd49}: color_data = 12'h4b3;
			{8'd148, 8'd50}: color_data = 12'h4b3;
			{8'd148, 8'd51}: color_data = 12'h4b3;
			{8'd148, 8'd52}: color_data = 12'h4b3;
			{8'd148, 8'd53}: color_data = 12'h4b3;
			{8'd148, 8'd54}: color_data = 12'h4b3;
			{8'd148, 8'd55}: color_data = 12'h4b3;
			{8'd148, 8'd56}: color_data = 12'h4a3;
			{8'd148, 8'd57}: color_data = 12'h4a3;
			{8'd148, 8'd58}: color_data = 12'h4a3;
			{8'd148, 8'd59}: color_data = 12'h4a3;
			{8'd148, 8'd60}: color_data = 12'h4a3;
			{8'd148, 8'd61}: color_data = 12'h4a3;
			{8'd148, 8'd62}: color_data = 12'h4a3;
			{8'd148, 8'd63}: color_data = 12'h4a3;
			{8'd148, 8'd64}: color_data = 12'h4a3;
			{8'd148, 8'd65}: color_data = 12'h4b3;
			{8'd148, 8'd66}: color_data = 12'h4a3;
			{8'd148, 8'd67}: color_data = 12'h020;
			{8'd148, 8'd68}: color_data = 12'h000;
			{8'd148, 8'd69}: color_data = 12'h000;
			{8'd148, 8'd70}: color_data = 12'h000;
			{8'd148, 8'd71}: color_data = 12'h000;
			{8'd148, 8'd72}: color_data = 12'h000;
			{8'd148, 8'd73}: color_data = 12'h000;
			{8'd148, 8'd74}: color_data = 12'h000;
			{8'd148, 8'd103}: color_data = 12'he00;
			{8'd148, 8'd104}: color_data = 12'he00;
			{8'd148, 8'd105}: color_data = 12'he00;
			{8'd148, 8'd106}: color_data = 12'he00;
			{8'd148, 8'd107}: color_data = 12'he00;
			{8'd148, 8'd108}: color_data = 12'he00;
			{8'd148, 8'd109}: color_data = 12'he01;
			{8'd148, 8'd110}: color_data = 12'he00;
			{8'd148, 8'd111}: color_data = 12'he01;
			{8'd148, 8'd133}: color_data = 12'he01;
			{8'd148, 8'd134}: color_data = 12'he00;
			{8'd148, 8'd135}: color_data = 12'he00;
			{8'd148, 8'd136}: color_data = 12'he00;
			{8'd148, 8'd137}: color_data = 12'he00;
			{8'd148, 8'd138}: color_data = 12'he00;
			{8'd148, 8'd139}: color_data = 12'he00;
			{8'd148, 8'd140}: color_data = 12'he00;
			{8'd148, 8'd141}: color_data = 12'he01;
			{8'd149, 8'd34}: color_data = 12'h000;
			{8'd149, 8'd35}: color_data = 12'h000;
			{8'd149, 8'd36}: color_data = 12'h000;
			{8'd149, 8'd37}: color_data = 12'h392;
			{8'd149, 8'd38}: color_data = 12'h4b3;
			{8'd149, 8'd39}: color_data = 12'h4a3;
			{8'd149, 8'd40}: color_data = 12'h4a3;
			{8'd149, 8'd41}: color_data = 12'h4a3;
			{8'd149, 8'd42}: color_data = 12'h4a3;
			{8'd149, 8'd43}: color_data = 12'h4a3;
			{8'd149, 8'd44}: color_data = 12'h4a3;
			{8'd149, 8'd45}: color_data = 12'h4a3;
			{8'd149, 8'd46}: color_data = 12'h4a3;
			{8'd149, 8'd47}: color_data = 12'h4a3;
			{8'd149, 8'd48}: color_data = 12'h4a3;
			{8'd149, 8'd49}: color_data = 12'h4a3;
			{8'd149, 8'd50}: color_data = 12'h4a3;
			{8'd149, 8'd51}: color_data = 12'h4a3;
			{8'd149, 8'd52}: color_data = 12'h4a3;
			{8'd149, 8'd53}: color_data = 12'h4a3;
			{8'd149, 8'd54}: color_data = 12'h4a3;
			{8'd149, 8'd55}: color_data = 12'h4a3;
			{8'd149, 8'd56}: color_data = 12'h4a3;
			{8'd149, 8'd57}: color_data = 12'h4a3;
			{8'd149, 8'd58}: color_data = 12'h4a3;
			{8'd149, 8'd59}: color_data = 12'h4a3;
			{8'd149, 8'd60}: color_data = 12'h4a3;
			{8'd149, 8'd61}: color_data = 12'h4a3;
			{8'd149, 8'd62}: color_data = 12'h4a3;
			{8'd149, 8'd63}: color_data = 12'h4a3;
			{8'd149, 8'd64}: color_data = 12'h4a3;
			{8'd149, 8'd65}: color_data = 12'h4b3;
			{8'd149, 8'd66}: color_data = 12'h372;
			{8'd149, 8'd67}: color_data = 12'h000;
			{8'd149, 8'd68}: color_data = 12'h000;
			{8'd149, 8'd69}: color_data = 12'h000;
			{8'd149, 8'd70}: color_data = 12'h000;
			{8'd149, 8'd71}: color_data = 12'h000;
			{8'd149, 8'd72}: color_data = 12'h000;
			{8'd149, 8'd73}: color_data = 12'h000;
			{8'd149, 8'd104}: color_data = 12'he00;
			{8'd149, 8'd105}: color_data = 12'he01;
			{8'd149, 8'd106}: color_data = 12'he00;
			{8'd149, 8'd107}: color_data = 12'he00;
			{8'd149, 8'd108}: color_data = 12'he00;
			{8'd149, 8'd109}: color_data = 12'he00;
			{8'd149, 8'd110}: color_data = 12'he00;
			{8'd149, 8'd111}: color_data = 12'he00;
			{8'd149, 8'd112}: color_data = 12'he00;
			{8'd149, 8'd132}: color_data = 12'he01;
			{8'd149, 8'd133}: color_data = 12'he00;
			{8'd149, 8'd134}: color_data = 12'he00;
			{8'd149, 8'd135}: color_data = 12'he00;
			{8'd149, 8'd136}: color_data = 12'he00;
			{8'd149, 8'd137}: color_data = 12'he00;
			{8'd149, 8'd138}: color_data = 12'he00;
			{8'd149, 8'd139}: color_data = 12'he00;
			{8'd149, 8'd140}: color_data = 12'he00;
			{8'd150, 8'd34}: color_data = 12'h000;
			{8'd150, 8'd35}: color_data = 12'h000;
			{8'd150, 8'd36}: color_data = 12'h000;
			{8'd150, 8'd37}: color_data = 12'h382;
			{8'd150, 8'd38}: color_data = 12'h4b3;
			{8'd150, 8'd39}: color_data = 12'h4a3;
			{8'd150, 8'd40}: color_data = 12'h4a3;
			{8'd150, 8'd41}: color_data = 12'h4a3;
			{8'd150, 8'd42}: color_data = 12'h4a3;
			{8'd150, 8'd43}: color_data = 12'h4a3;
			{8'd150, 8'd44}: color_data = 12'h4a3;
			{8'd150, 8'd45}: color_data = 12'h4a3;
			{8'd150, 8'd46}: color_data = 12'h4a3;
			{8'd150, 8'd47}: color_data = 12'h4a3;
			{8'd150, 8'd48}: color_data = 12'h4a3;
			{8'd150, 8'd49}: color_data = 12'h4a3;
			{8'd150, 8'd50}: color_data = 12'h4a3;
			{8'd150, 8'd51}: color_data = 12'h4a3;
			{8'd150, 8'd52}: color_data = 12'h4a3;
			{8'd150, 8'd53}: color_data = 12'h4a3;
			{8'd150, 8'd54}: color_data = 12'h4a3;
			{8'd150, 8'd55}: color_data = 12'h4a3;
			{8'd150, 8'd56}: color_data = 12'h4a3;
			{8'd150, 8'd57}: color_data = 12'h4a3;
			{8'd150, 8'd58}: color_data = 12'h4a3;
			{8'd150, 8'd59}: color_data = 12'h4a3;
			{8'd150, 8'd60}: color_data = 12'h4a3;
			{8'd150, 8'd61}: color_data = 12'h4a3;
			{8'd150, 8'd62}: color_data = 12'h4a3;
			{8'd150, 8'd63}: color_data = 12'h4a3;
			{8'd150, 8'd64}: color_data = 12'h4b3;
			{8'd150, 8'd65}: color_data = 12'h4b3;
			{8'd150, 8'd66}: color_data = 12'h131;
			{8'd150, 8'd67}: color_data = 12'h000;
			{8'd150, 8'd68}: color_data = 12'h000;
			{8'd150, 8'd69}: color_data = 12'h000;
			{8'd150, 8'd70}: color_data = 12'h000;
			{8'd150, 8'd71}: color_data = 12'h000;
			{8'd150, 8'd72}: color_data = 12'h000;
			{8'd150, 8'd73}: color_data = 12'h000;
			{8'd150, 8'd104}: color_data = 12'hc00;
			{8'd150, 8'd105}: color_data = 12'he00;
			{8'd150, 8'd106}: color_data = 12'hf01;
			{8'd150, 8'd107}: color_data = 12'he00;
			{8'd150, 8'd108}: color_data = 12'he00;
			{8'd150, 8'd109}: color_data = 12'he00;
			{8'd150, 8'd110}: color_data = 12'he00;
			{8'd150, 8'd111}: color_data = 12'he01;
			{8'd150, 8'd112}: color_data = 12'he00;
			{8'd150, 8'd113}: color_data = 12'he00;
			{8'd150, 8'd130}: color_data = 12'hc00;
			{8'd150, 8'd131}: color_data = 12'he00;
			{8'd150, 8'd132}: color_data = 12'he00;
			{8'd150, 8'd133}: color_data = 12'he00;
			{8'd150, 8'd134}: color_data = 12'he00;
			{8'd150, 8'd135}: color_data = 12'he00;
			{8'd150, 8'd136}: color_data = 12'he00;
			{8'd150, 8'd137}: color_data = 12'he00;
			{8'd150, 8'd138}: color_data = 12'hf01;
			{8'd150, 8'd139}: color_data = 12'he00;
			{8'd151, 8'd34}: color_data = 12'h000;
			{8'd151, 8'd35}: color_data = 12'h000;
			{8'd151, 8'd36}: color_data = 12'h000;
			{8'd151, 8'd37}: color_data = 12'h120;
			{8'd151, 8'd38}: color_data = 12'h393;
			{8'd151, 8'd39}: color_data = 12'h4b3;
			{8'd151, 8'd40}: color_data = 12'h4a3;
			{8'd151, 8'd41}: color_data = 12'h4a3;
			{8'd151, 8'd42}: color_data = 12'h4a3;
			{8'd151, 8'd43}: color_data = 12'h4a3;
			{8'd151, 8'd44}: color_data = 12'h4a3;
			{8'd151, 8'd45}: color_data = 12'h4a3;
			{8'd151, 8'd46}: color_data = 12'h4a3;
			{8'd151, 8'd47}: color_data = 12'h4a3;
			{8'd151, 8'd48}: color_data = 12'h4a3;
			{8'd151, 8'd49}: color_data = 12'h4a3;
			{8'd151, 8'd50}: color_data = 12'h4a3;
			{8'd151, 8'd51}: color_data = 12'h4a3;
			{8'd151, 8'd52}: color_data = 12'h4a3;
			{8'd151, 8'd53}: color_data = 12'h4a3;
			{8'd151, 8'd54}: color_data = 12'h4a3;
			{8'd151, 8'd55}: color_data = 12'h4a3;
			{8'd151, 8'd56}: color_data = 12'h4a3;
			{8'd151, 8'd57}: color_data = 12'h4a3;
			{8'd151, 8'd58}: color_data = 12'h4a3;
			{8'd151, 8'd59}: color_data = 12'h4a3;
			{8'd151, 8'd60}: color_data = 12'h4a3;
			{8'd151, 8'd61}: color_data = 12'h4a3;
			{8'd151, 8'd62}: color_data = 12'h4a3;
			{8'd151, 8'd63}: color_data = 12'h4a3;
			{8'd151, 8'd64}: color_data = 12'h4b3;
			{8'd151, 8'd65}: color_data = 12'h382;
			{8'd151, 8'd66}: color_data = 12'h000;
			{8'd151, 8'd67}: color_data = 12'h000;
			{8'd151, 8'd68}: color_data = 12'h000;
			{8'd151, 8'd69}: color_data = 12'h000;
			{8'd151, 8'd70}: color_data = 12'h000;
			{8'd151, 8'd71}: color_data = 12'h000;
			{8'd151, 8'd72}: color_data = 12'h000;
			{8'd151, 8'd73}: color_data = 12'h000;
			{8'd151, 8'd105}: color_data = 12'he00;
			{8'd151, 8'd106}: color_data = 12'he00;
			{8'd151, 8'd107}: color_data = 12'hf01;
			{8'd151, 8'd108}: color_data = 12'he00;
			{8'd151, 8'd109}: color_data = 12'he00;
			{8'd151, 8'd110}: color_data = 12'he00;
			{8'd151, 8'd111}: color_data = 12'he00;
			{8'd151, 8'd112}: color_data = 12'he00;
			{8'd151, 8'd113}: color_data = 12'he00;
			{8'd151, 8'd114}: color_data = 12'he00;
			{8'd151, 8'd115}: color_data = 12'he00;
			{8'd151, 8'd116}: color_data = 12'hf00;
			{8'd151, 8'd128}: color_data = 12'hc00;
			{8'd151, 8'd129}: color_data = 12'he00;
			{8'd151, 8'd130}: color_data = 12'he00;
			{8'd151, 8'd131}: color_data = 12'he01;
			{8'd151, 8'd132}: color_data = 12'he00;
			{8'd151, 8'd133}: color_data = 12'he00;
			{8'd151, 8'd134}: color_data = 12'he00;
			{8'd151, 8'd135}: color_data = 12'he00;
			{8'd151, 8'd136}: color_data = 12'he00;
			{8'd151, 8'd137}: color_data = 12'hf01;
			{8'd151, 8'd138}: color_data = 12'he00;
			{8'd151, 8'd139}: color_data = 12'hd00;
			{8'd152, 8'd34}: color_data = 12'h000;
			{8'd152, 8'd35}: color_data = 12'h000;
			{8'd152, 8'd36}: color_data = 12'h000;
			{8'd152, 8'd37}: color_data = 12'h000;
			{8'd152, 8'd38}: color_data = 12'h010;
			{8'd152, 8'd39}: color_data = 12'h272;
			{8'd152, 8'd40}: color_data = 12'h4b3;
			{8'd152, 8'd41}: color_data = 12'h4b3;
			{8'd152, 8'd42}: color_data = 12'h4a3;
			{8'd152, 8'd43}: color_data = 12'h4a3;
			{8'd152, 8'd44}: color_data = 12'h4a3;
			{8'd152, 8'd45}: color_data = 12'h4a3;
			{8'd152, 8'd46}: color_data = 12'h4a3;
			{8'd152, 8'd47}: color_data = 12'h4a3;
			{8'd152, 8'd48}: color_data = 12'h4a3;
			{8'd152, 8'd49}: color_data = 12'h4a3;
			{8'd152, 8'd50}: color_data = 12'h4a3;
			{8'd152, 8'd51}: color_data = 12'h4a3;
			{8'd152, 8'd52}: color_data = 12'h4a3;
			{8'd152, 8'd53}: color_data = 12'h4a3;
			{8'd152, 8'd54}: color_data = 12'h4a3;
			{8'd152, 8'd55}: color_data = 12'h4a3;
			{8'd152, 8'd56}: color_data = 12'h4a3;
			{8'd152, 8'd57}: color_data = 12'h4a3;
			{8'd152, 8'd58}: color_data = 12'h4a3;
			{8'd152, 8'd59}: color_data = 12'h4a3;
			{8'd152, 8'd60}: color_data = 12'h4a3;
			{8'd152, 8'd61}: color_data = 12'h4a3;
			{8'd152, 8'd62}: color_data = 12'h4a3;
			{8'd152, 8'd63}: color_data = 12'h4a3;
			{8'd152, 8'd64}: color_data = 12'h4b3;
			{8'd152, 8'd65}: color_data = 12'h141;
			{8'd152, 8'd66}: color_data = 12'h000;
			{8'd152, 8'd67}: color_data = 12'h000;
			{8'd152, 8'd68}: color_data = 12'h000;
			{8'd152, 8'd69}: color_data = 12'h000;
			{8'd152, 8'd70}: color_data = 12'h000;
			{8'd152, 8'd71}: color_data = 12'h000;
			{8'd152, 8'd72}: color_data = 12'h000;
			{8'd152, 8'd106}: color_data = 12'he01;
			{8'd152, 8'd107}: color_data = 12'he00;
			{8'd152, 8'd108}: color_data = 12'he01;
			{8'd152, 8'd109}: color_data = 12'he00;
			{8'd152, 8'd110}: color_data = 12'he00;
			{8'd152, 8'd111}: color_data = 12'he00;
			{8'd152, 8'd112}: color_data = 12'he00;
			{8'd152, 8'd113}: color_data = 12'he00;
			{8'd152, 8'd114}: color_data = 12'he01;
			{8'd152, 8'd115}: color_data = 12'he00;
			{8'd152, 8'd116}: color_data = 12'he00;
			{8'd152, 8'd117}: color_data = 12'he00;
			{8'd152, 8'd118}: color_data = 12'he01;
			{8'd152, 8'd119}: color_data = 12'hd01;
			{8'd152, 8'd124}: color_data = 12'hf00;
			{8'd152, 8'd125}: color_data = 12'hd00;
			{8'd152, 8'd126}: color_data = 12'he00;
			{8'd152, 8'd127}: color_data = 12'he00;
			{8'd152, 8'd128}: color_data = 12'he00;
			{8'd152, 8'd129}: color_data = 12'he01;
			{8'd152, 8'd130}: color_data = 12'he01;
			{8'd152, 8'd131}: color_data = 12'he00;
			{8'd152, 8'd132}: color_data = 12'he00;
			{8'd152, 8'd133}: color_data = 12'he00;
			{8'd152, 8'd134}: color_data = 12'he00;
			{8'd152, 8'd135}: color_data = 12'he00;
			{8'd152, 8'd136}: color_data = 12'hf01;
			{8'd152, 8'd137}: color_data = 12'he00;
			{8'd152, 8'd138}: color_data = 12'he01;
			{8'd153, 8'd35}: color_data = 12'h000;
			{8'd153, 8'd36}: color_data = 12'h000;
			{8'd153, 8'd37}: color_data = 12'h000;
			{8'd153, 8'd38}: color_data = 12'h000;
			{8'd153, 8'd39}: color_data = 12'h000;
			{8'd153, 8'd40}: color_data = 12'h141;
			{8'd153, 8'd41}: color_data = 12'h4a3;
			{8'd153, 8'd42}: color_data = 12'h4b3;
			{8'd153, 8'd43}: color_data = 12'h4a3;
			{8'd153, 8'd44}: color_data = 12'h4a3;
			{8'd153, 8'd45}: color_data = 12'h4a3;
			{8'd153, 8'd46}: color_data = 12'h4a3;
			{8'd153, 8'd47}: color_data = 12'h4a3;
			{8'd153, 8'd48}: color_data = 12'h4a3;
			{8'd153, 8'd49}: color_data = 12'h4a3;
			{8'd153, 8'd50}: color_data = 12'h4a3;
			{8'd153, 8'd51}: color_data = 12'h4a3;
			{8'd153, 8'd52}: color_data = 12'h4a3;
			{8'd153, 8'd53}: color_data = 12'h4a3;
			{8'd153, 8'd54}: color_data = 12'h4a3;
			{8'd153, 8'd55}: color_data = 12'h4a3;
			{8'd153, 8'd56}: color_data = 12'h4a3;
			{8'd153, 8'd57}: color_data = 12'h4a3;
			{8'd153, 8'd58}: color_data = 12'h4a3;
			{8'd153, 8'd59}: color_data = 12'h4a3;
			{8'd153, 8'd60}: color_data = 12'h4a3;
			{8'd153, 8'd61}: color_data = 12'h4a3;
			{8'd153, 8'd62}: color_data = 12'h4a3;
			{8'd153, 8'd63}: color_data = 12'h4b3;
			{8'd153, 8'd64}: color_data = 12'h392;
			{8'd153, 8'd65}: color_data = 12'h000;
			{8'd153, 8'd66}: color_data = 12'h000;
			{8'd153, 8'd67}: color_data = 12'h000;
			{8'd153, 8'd68}: color_data = 12'h000;
			{8'd153, 8'd69}: color_data = 12'h000;
			{8'd153, 8'd70}: color_data = 12'h000;
			{8'd153, 8'd71}: color_data = 12'h000;
			{8'd153, 8'd72}: color_data = 12'h000;
			{8'd153, 8'd107}: color_data = 12'hd00;
			{8'd153, 8'd108}: color_data = 12'he00;
			{8'd153, 8'd109}: color_data = 12'hf01;
			{8'd153, 8'd110}: color_data = 12'he00;
			{8'd153, 8'd111}: color_data = 12'he00;
			{8'd153, 8'd112}: color_data = 12'he00;
			{8'd153, 8'd113}: color_data = 12'he00;
			{8'd153, 8'd114}: color_data = 12'he00;
			{8'd153, 8'd115}: color_data = 12'he00;
			{8'd153, 8'd116}: color_data = 12'he00;
			{8'd153, 8'd117}: color_data = 12'he01;
			{8'd153, 8'd118}: color_data = 12'he00;
			{8'd153, 8'd119}: color_data = 12'he00;
			{8'd153, 8'd120}: color_data = 12'he00;
			{8'd153, 8'd121}: color_data = 12'he00;
			{8'd153, 8'd122}: color_data = 12'he00;
			{8'd153, 8'd123}: color_data = 12'he00;
			{8'd153, 8'd124}: color_data = 12'he00;
			{8'd153, 8'd125}: color_data = 12'he00;
			{8'd153, 8'd126}: color_data = 12'he00;
			{8'd153, 8'd127}: color_data = 12'he01;
			{8'd153, 8'd128}: color_data = 12'he00;
			{8'd153, 8'd129}: color_data = 12'he00;
			{8'd153, 8'd130}: color_data = 12'he00;
			{8'd153, 8'd131}: color_data = 12'he00;
			{8'd153, 8'd132}: color_data = 12'he00;
			{8'd153, 8'd133}: color_data = 12'he00;
			{8'd153, 8'd134}: color_data = 12'he00;
			{8'd153, 8'd135}: color_data = 12'he01;
			{8'd153, 8'd136}: color_data = 12'he00;
			{8'd153, 8'd137}: color_data = 12'he00;
			{8'd154, 8'd36}: color_data = 12'h000;
			{8'd154, 8'd37}: color_data = 12'h000;
			{8'd154, 8'd38}: color_data = 12'h000;
			{8'd154, 8'd39}: color_data = 12'h000;
			{8'd154, 8'd40}: color_data = 12'h000;
			{8'd154, 8'd41}: color_data = 12'h020;
			{8'd154, 8'd42}: color_data = 12'h382;
			{8'd154, 8'd43}: color_data = 12'h4b3;
			{8'd154, 8'd44}: color_data = 12'h4b3;
			{8'd154, 8'd45}: color_data = 12'h4a3;
			{8'd154, 8'd46}: color_data = 12'h4a3;
			{8'd154, 8'd47}: color_data = 12'h4a3;
			{8'd154, 8'd48}: color_data = 12'h4a3;
			{8'd154, 8'd49}: color_data = 12'h4a3;
			{8'd154, 8'd50}: color_data = 12'h4a3;
			{8'd154, 8'd51}: color_data = 12'h4a3;
			{8'd154, 8'd52}: color_data = 12'h4a3;
			{8'd154, 8'd53}: color_data = 12'h4a3;
			{8'd154, 8'd54}: color_data = 12'h4a3;
			{8'd154, 8'd55}: color_data = 12'h4a3;
			{8'd154, 8'd56}: color_data = 12'h4a3;
			{8'd154, 8'd57}: color_data = 12'h4a3;
			{8'd154, 8'd58}: color_data = 12'h4a3;
			{8'd154, 8'd59}: color_data = 12'h4a3;
			{8'd154, 8'd60}: color_data = 12'h4a3;
			{8'd154, 8'd61}: color_data = 12'h4a3;
			{8'd154, 8'd62}: color_data = 12'h4a3;
			{8'd154, 8'd63}: color_data = 12'h4b3;
			{8'd154, 8'd64}: color_data = 12'h151;
			{8'd154, 8'd65}: color_data = 12'h000;
			{8'd154, 8'd66}: color_data = 12'h000;
			{8'd154, 8'd67}: color_data = 12'h000;
			{8'd154, 8'd68}: color_data = 12'h000;
			{8'd154, 8'd69}: color_data = 12'h000;
			{8'd154, 8'd70}: color_data = 12'h000;
			{8'd154, 8'd71}: color_data = 12'h000;
			{8'd154, 8'd108}: color_data = 12'he01;
			{8'd154, 8'd109}: color_data = 12'he00;
			{8'd154, 8'd110}: color_data = 12'he00;
			{8'd154, 8'd111}: color_data = 12'he00;
			{8'd154, 8'd112}: color_data = 12'he00;
			{8'd154, 8'd113}: color_data = 12'he00;
			{8'd154, 8'd114}: color_data = 12'he00;
			{8'd154, 8'd115}: color_data = 12'he00;
			{8'd154, 8'd116}: color_data = 12'he00;
			{8'd154, 8'd117}: color_data = 12'he00;
			{8'd154, 8'd118}: color_data = 12'he00;
			{8'd154, 8'd119}: color_data = 12'he00;
			{8'd154, 8'd120}: color_data = 12'he00;
			{8'd154, 8'd121}: color_data = 12'he00;
			{8'd154, 8'd122}: color_data = 12'he01;
			{8'd154, 8'd123}: color_data = 12'he00;
			{8'd154, 8'd124}: color_data = 12'he00;
			{8'd154, 8'd125}: color_data = 12'he00;
			{8'd154, 8'd126}: color_data = 12'he00;
			{8'd154, 8'd127}: color_data = 12'he00;
			{8'd154, 8'd128}: color_data = 12'he00;
			{8'd154, 8'd129}: color_data = 12'he00;
			{8'd154, 8'd130}: color_data = 12'he00;
			{8'd154, 8'd131}: color_data = 12'he00;
			{8'd154, 8'd132}: color_data = 12'he00;
			{8'd154, 8'd133}: color_data = 12'he01;
			{8'd154, 8'd134}: color_data = 12'he00;
			{8'd154, 8'd135}: color_data = 12'he01;
			{8'd154, 8'd136}: color_data = 12'hf00;
			{8'd155, 8'd38}: color_data = 12'h000;
			{8'd155, 8'd39}: color_data = 12'h000;
			{8'd155, 8'd40}: color_data = 12'h000;
			{8'd155, 8'd41}: color_data = 12'h000;
			{8'd155, 8'd42}: color_data = 12'h000;
			{8'd155, 8'd43}: color_data = 12'h251;
			{8'd155, 8'd44}: color_data = 12'h4a3;
			{8'd155, 8'd45}: color_data = 12'h4b3;
			{8'd155, 8'd46}: color_data = 12'h4a3;
			{8'd155, 8'd47}: color_data = 12'h4a3;
			{8'd155, 8'd48}: color_data = 12'h4a3;
			{8'd155, 8'd49}: color_data = 12'h4a3;
			{8'd155, 8'd50}: color_data = 12'h4a3;
			{8'd155, 8'd51}: color_data = 12'h4a3;
			{8'd155, 8'd52}: color_data = 12'h4a3;
			{8'd155, 8'd53}: color_data = 12'h4a3;
			{8'd155, 8'd54}: color_data = 12'h4a3;
			{8'd155, 8'd55}: color_data = 12'h4a3;
			{8'd155, 8'd56}: color_data = 12'h4a3;
			{8'd155, 8'd57}: color_data = 12'h4a3;
			{8'd155, 8'd58}: color_data = 12'h4a3;
			{8'd155, 8'd59}: color_data = 12'h4b3;
			{8'd155, 8'd60}: color_data = 12'h4b3;
			{8'd155, 8'd61}: color_data = 12'h4b3;
			{8'd155, 8'd62}: color_data = 12'h4b3;
			{8'd155, 8'd63}: color_data = 12'h392;
			{8'd155, 8'd64}: color_data = 12'h010;
			{8'd155, 8'd65}: color_data = 12'h000;
			{8'd155, 8'd66}: color_data = 12'h000;
			{8'd155, 8'd67}: color_data = 12'h000;
			{8'd155, 8'd68}: color_data = 12'h000;
			{8'd155, 8'd69}: color_data = 12'h000;
			{8'd155, 8'd70}: color_data = 12'h000;
			{8'd155, 8'd71}: color_data = 12'h000;
			{8'd155, 8'd110}: color_data = 12'he00;
			{8'd155, 8'd111}: color_data = 12'he00;
			{8'd155, 8'd112}: color_data = 12'he01;
			{8'd155, 8'd113}: color_data = 12'he00;
			{8'd155, 8'd114}: color_data = 12'he00;
			{8'd155, 8'd115}: color_data = 12'he00;
			{8'd155, 8'd116}: color_data = 12'he00;
			{8'd155, 8'd117}: color_data = 12'he00;
			{8'd155, 8'd118}: color_data = 12'he00;
			{8'd155, 8'd119}: color_data = 12'he00;
			{8'd155, 8'd120}: color_data = 12'he00;
			{8'd155, 8'd121}: color_data = 12'he00;
			{8'd155, 8'd122}: color_data = 12'he00;
			{8'd155, 8'd123}: color_data = 12'he00;
			{8'd155, 8'd124}: color_data = 12'he00;
			{8'd155, 8'd125}: color_data = 12'he00;
			{8'd155, 8'd126}: color_data = 12'he00;
			{8'd155, 8'd127}: color_data = 12'he00;
			{8'd155, 8'd128}: color_data = 12'he00;
			{8'd155, 8'd129}: color_data = 12'he00;
			{8'd155, 8'd130}: color_data = 12'he00;
			{8'd155, 8'd131}: color_data = 12'he00;
			{8'd155, 8'd132}: color_data = 12'he00;
			{8'd155, 8'd133}: color_data = 12'he00;
			{8'd155, 8'd134}: color_data = 12'he00;
			{8'd156, 8'd39}: color_data = 12'h000;
			{8'd156, 8'd40}: color_data = 12'h000;
			{8'd156, 8'd41}: color_data = 12'h000;
			{8'd156, 8'd42}: color_data = 12'h000;
			{8'd156, 8'd43}: color_data = 12'h000;
			{8'd156, 8'd44}: color_data = 12'h130;
			{8'd156, 8'd45}: color_data = 12'h392;
			{8'd156, 8'd46}: color_data = 12'h4b3;
			{8'd156, 8'd47}: color_data = 12'h4a3;
			{8'd156, 8'd48}: color_data = 12'h4a3;
			{8'd156, 8'd49}: color_data = 12'h4a3;
			{8'd156, 8'd50}: color_data = 12'h4a3;
			{8'd156, 8'd51}: color_data = 12'h4a3;
			{8'd156, 8'd52}: color_data = 12'h4a3;
			{8'd156, 8'd53}: color_data = 12'h4a3;
			{8'd156, 8'd54}: color_data = 12'h4a3;
			{8'd156, 8'd55}: color_data = 12'h4a3;
			{8'd156, 8'd56}: color_data = 12'h4b3;
			{8'd156, 8'd57}: color_data = 12'h4b3;
			{8'd156, 8'd58}: color_data = 12'h4b3;
			{8'd156, 8'd59}: color_data = 12'h4b3;
			{8'd156, 8'd60}: color_data = 12'h392;
			{8'd156, 8'd61}: color_data = 12'h272;
			{8'd156, 8'd62}: color_data = 12'h151;
			{8'd156, 8'd63}: color_data = 12'h010;
			{8'd156, 8'd64}: color_data = 12'h000;
			{8'd156, 8'd65}: color_data = 12'h000;
			{8'd156, 8'd66}: color_data = 12'h000;
			{8'd156, 8'd67}: color_data = 12'h000;
			{8'd156, 8'd68}: color_data = 12'h000;
			{8'd156, 8'd69}: color_data = 12'h000;
			{8'd156, 8'd70}: color_data = 12'h000;
			{8'd156, 8'd111}: color_data = 12'he01;
			{8'd156, 8'd112}: color_data = 12'he00;
			{8'd156, 8'd113}: color_data = 12'he00;
			{8'd156, 8'd114}: color_data = 12'he01;
			{8'd156, 8'd115}: color_data = 12'he01;
			{8'd156, 8'd116}: color_data = 12'he00;
			{8'd156, 8'd117}: color_data = 12'he00;
			{8'd156, 8'd118}: color_data = 12'he00;
			{8'd156, 8'd119}: color_data = 12'he00;
			{8'd156, 8'd120}: color_data = 12'he00;
			{8'd156, 8'd121}: color_data = 12'he00;
			{8'd156, 8'd122}: color_data = 12'he00;
			{8'd156, 8'd123}: color_data = 12'he00;
			{8'd156, 8'd124}: color_data = 12'he00;
			{8'd156, 8'd125}: color_data = 12'he00;
			{8'd156, 8'd126}: color_data = 12'he00;
			{8'd156, 8'd127}: color_data = 12'he00;
			{8'd156, 8'd128}: color_data = 12'he00;
			{8'd156, 8'd129}: color_data = 12'he01;
			{8'd156, 8'd130}: color_data = 12'he00;
			{8'd156, 8'd131}: color_data = 12'he00;
			{8'd156, 8'd132}: color_data = 12'he00;
			{8'd156, 8'd133}: color_data = 12'hf00;
			{8'd157, 8'd40}: color_data = 12'h000;
			{8'd157, 8'd41}: color_data = 12'h000;
			{8'd157, 8'd42}: color_data = 12'h000;
			{8'd157, 8'd43}: color_data = 12'h000;
			{8'd157, 8'd44}: color_data = 12'h000;
			{8'd157, 8'd45}: color_data = 12'h010;
			{8'd157, 8'd46}: color_data = 12'h272;
			{8'd157, 8'd47}: color_data = 12'h4b3;
			{8'd157, 8'd48}: color_data = 12'h4b3;
			{8'd157, 8'd49}: color_data = 12'h4a3;
			{8'd157, 8'd50}: color_data = 12'h4a3;
			{8'd157, 8'd51}: color_data = 12'h4a3;
			{8'd157, 8'd52}: color_data = 12'h4b3;
			{8'd157, 8'd53}: color_data = 12'h4b3;
			{8'd157, 8'd54}: color_data = 12'h4b3;
			{8'd157, 8'd55}: color_data = 12'h4b3;
			{8'd157, 8'd56}: color_data = 12'h393;
			{8'd157, 8'd57}: color_data = 12'h372;
			{8'd157, 8'd58}: color_data = 12'h251;
			{8'd157, 8'd59}: color_data = 12'h120;
			{8'd157, 8'd60}: color_data = 12'h000;
			{8'd157, 8'd61}: color_data = 12'h000;
			{8'd157, 8'd62}: color_data = 12'h000;
			{8'd157, 8'd63}: color_data = 12'h000;
			{8'd157, 8'd64}: color_data = 12'h000;
			{8'd157, 8'd65}: color_data = 12'h000;
			{8'd157, 8'd66}: color_data = 12'h000;
			{8'd157, 8'd67}: color_data = 12'h000;
			{8'd157, 8'd68}: color_data = 12'h000;
			{8'd157, 8'd69}: color_data = 12'h000;
			{8'd157, 8'd70}: color_data = 12'h000;
			{8'd157, 8'd113}: color_data = 12'he01;
			{8'd157, 8'd114}: color_data = 12'he00;
			{8'd157, 8'd115}: color_data = 12'he00;
			{8'd157, 8'd116}: color_data = 12'he00;
			{8'd157, 8'd117}: color_data = 12'he00;
			{8'd157, 8'd118}: color_data = 12'he01;
			{8'd157, 8'd119}: color_data = 12'he01;
			{8'd157, 8'd120}: color_data = 12'he01;
			{8'd157, 8'd121}: color_data = 12'he00;
			{8'd157, 8'd122}: color_data = 12'he00;
			{8'd157, 8'd123}: color_data = 12'he00;
			{8'd157, 8'd124}: color_data = 12'he01;
			{8'd157, 8'd125}: color_data = 12'he01;
			{8'd157, 8'd126}: color_data = 12'he01;
			{8'd157, 8'd127}: color_data = 12'he00;
			{8'd157, 8'd128}: color_data = 12'he00;
			{8'd157, 8'd129}: color_data = 12'he00;
			{8'd157, 8'd130}: color_data = 12'he00;
			{8'd157, 8'd131}: color_data = 12'hc00;
			{8'd158, 8'd42}: color_data = 12'h000;
			{8'd158, 8'd43}: color_data = 12'h000;
			{8'd158, 8'd44}: color_data = 12'h000;
			{8'd158, 8'd45}: color_data = 12'h000;
			{8'd158, 8'd46}: color_data = 12'h000;
			{8'd158, 8'd47}: color_data = 12'h141;
			{8'd158, 8'd48}: color_data = 12'h4a3;
			{8'd158, 8'd49}: color_data = 12'h4b3;
			{8'd158, 8'd50}: color_data = 12'h4b3;
			{8'd158, 8'd51}: color_data = 12'h4b3;
			{8'd158, 8'd52}: color_data = 12'h393;
			{8'd158, 8'd53}: color_data = 12'h372;
			{8'd158, 8'd54}: color_data = 12'h251;
			{8'd158, 8'd55}: color_data = 12'h120;
			{8'd158, 8'd56}: color_data = 12'h000;
			{8'd158, 8'd57}: color_data = 12'h000;
			{8'd158, 8'd58}: color_data = 12'h000;
			{8'd158, 8'd59}: color_data = 12'h000;
			{8'd158, 8'd60}: color_data = 12'h000;
			{8'd158, 8'd61}: color_data = 12'h000;
			{8'd158, 8'd62}: color_data = 12'h000;
			{8'd158, 8'd63}: color_data = 12'h000;
			{8'd158, 8'd64}: color_data = 12'h000;
			{8'd158, 8'd65}: color_data = 12'h000;
			{8'd158, 8'd66}: color_data = 12'h000;
			{8'd158, 8'd67}: color_data = 12'h000;
			{8'd158, 8'd68}: color_data = 12'h000;
			{8'd158, 8'd69}: color_data = 12'h000;
			{8'd158, 8'd116}: color_data = 12'he01;
			{8'd158, 8'd117}: color_data = 12'he00;
			{8'd158, 8'd118}: color_data = 12'he00;
			{8'd158, 8'd119}: color_data = 12'he00;
			{8'd158, 8'd120}: color_data = 12'he00;
			{8'd158, 8'd121}: color_data = 12'he00;
			{8'd158, 8'd122}: color_data = 12'he00;
			{8'd158, 8'd123}: color_data = 12'he00;
			{8'd158, 8'd124}: color_data = 12'he00;
			{8'd158, 8'd125}: color_data = 12'he00;
			{8'd158, 8'd126}: color_data = 12'he00;
			{8'd158, 8'd127}: color_data = 12'he00;
			{8'd158, 8'd128}: color_data = 12'he00;
			{8'd159, 8'd43}: color_data = 12'h000;
			{8'd159, 8'd44}: color_data = 12'h000;
			{8'd159, 8'd45}: color_data = 12'h000;
			{8'd159, 8'd46}: color_data = 12'h000;
			{8'd159, 8'd47}: color_data = 12'h000;
			{8'd159, 8'd48}: color_data = 12'h010;
			{8'd159, 8'd49}: color_data = 12'h262;
			{8'd159, 8'd50}: color_data = 12'h251;
			{8'd159, 8'd51}: color_data = 12'h120;
			{8'd159, 8'd52}: color_data = 12'h000;
			{8'd159, 8'd53}: color_data = 12'h000;
			{8'd159, 8'd54}: color_data = 12'h000;
			{8'd159, 8'd55}: color_data = 12'h000;
			{8'd159, 8'd56}: color_data = 12'h000;
			{8'd159, 8'd57}: color_data = 12'h000;
			{8'd159, 8'd58}: color_data = 12'h000;
			{8'd159, 8'd59}: color_data = 12'h000;
			{8'd159, 8'd60}: color_data = 12'h000;
			{8'd159, 8'd61}: color_data = 12'h000;
			{8'd159, 8'd62}: color_data = 12'h000;
			{8'd159, 8'd63}: color_data = 12'h000;
			{8'd159, 8'd64}: color_data = 12'h000;
			{8'd159, 8'd65}: color_data = 12'h000;
			{8'd159, 8'd66}: color_data = 12'h000;
			{8'd159, 8'd67}: color_data = 12'h000;
			{8'd160, 8'd45}: color_data = 12'h000;
			{8'd160, 8'd46}: color_data = 12'h000;
			{8'd160, 8'd47}: color_data = 12'h000;
			{8'd160, 8'd48}: color_data = 12'h000;
			{8'd160, 8'd49}: color_data = 12'h000;
			{8'd160, 8'd50}: color_data = 12'h000;
			{8'd160, 8'd51}: color_data = 12'h000;
			{8'd160, 8'd52}: color_data = 12'h000;
			{8'd160, 8'd53}: color_data = 12'h000;
			{8'd160, 8'd54}: color_data = 12'h000;
			{8'd160, 8'd55}: color_data = 12'h000;
			{8'd160, 8'd56}: color_data = 12'h000;
			{8'd160, 8'd57}: color_data = 12'h000;
			{8'd160, 8'd58}: color_data = 12'h000;
			{8'd160, 8'd59}: color_data = 12'h000;
			{8'd160, 8'd60}: color_data = 12'h000;
			{8'd160, 8'd61}: color_data = 12'h000;
			{8'd160, 8'd62}: color_data = 12'h000;
			{8'd160, 8'd63}: color_data = 12'h000;
			{8'd161, 8'd46}: color_data = 12'h000;
			{8'd161, 8'd47}: color_data = 12'h000;
			{8'd161, 8'd48}: color_data = 12'h000;
			{8'd161, 8'd49}: color_data = 12'h000;
			{8'd161, 8'd50}: color_data = 12'h000;
			{8'd161, 8'd51}: color_data = 12'h000;
			{8'd161, 8'd52}: color_data = 12'h000;
			{8'd161, 8'd53}: color_data = 12'h000;
			{8'd161, 8'd54}: color_data = 12'h000;
			{8'd161, 8'd55}: color_data = 12'h000;
			{8'd161, 8'd56}: color_data = 12'h000;
			{8'd161, 8'd57}: color_data = 12'h000;
			{8'd161, 8'd58}: color_data = 12'h000;
			{8'd161, 8'd59}: color_data = 12'h000;
			{8'd161, 8'd67}: color_data = 12'h000;
			{8'd161, 8'd68}: color_data = 12'h000;
			{8'd162, 8'd47}: color_data = 12'h000;
			{8'd162, 8'd48}: color_data = 12'h000;
			{8'd162, 8'd49}: color_data = 12'h000;
			{8'd162, 8'd50}: color_data = 12'h000;
			{8'd162, 8'd51}: color_data = 12'h000;
			{8'd162, 8'd52}: color_data = 12'h000;
			{8'd162, 8'd53}: color_data = 12'h000;
			{8'd162, 8'd54}: color_data = 12'h000;
			{8'd162, 8'd55}: color_data = 12'h000;
			{8'd162, 8'd67}: color_data = 12'h000;
			{8'd162, 8'd68}: color_data = 12'h000;
			{8'd162, 8'd69}: color_data = 12'h000;
			{8'd162, 8'd70}: color_data = 12'h000;
			{8'd162, 8'd71}: color_data = 12'h000;
			{8'd162, 8'd72}: color_data = 12'h000;
			{8'd163, 8'd67}: color_data = 12'h000;
			{8'd163, 8'd68}: color_data = 12'h000;
			{8'd163, 8'd69}: color_data = 12'h000;
			{8'd163, 8'd70}: color_data = 12'h000;
			{8'd163, 8'd71}: color_data = 12'h000;
			{8'd163, 8'd72}: color_data = 12'h000;
			{8'd164, 8'd67}: color_data = 12'h000;
			{8'd164, 8'd68}: color_data = 12'h000;
			{8'd164, 8'd70}: color_data = 12'h000;
			{8'd164, 8'd71}: color_data = 12'h000;
			{8'd164, 8'd72}: color_data = 12'h000;
			{8'd165, 8'd67}: color_data = 12'h000;
			{8'd165, 8'd68}: color_data = 12'h000;
			{8'd165, 8'd69}: color_data = 12'h000;
			{8'd165, 8'd70}: color_data = 12'h000;
			{8'd165, 8'd71}: color_data = 12'h000;
			{8'd165, 8'd72}: color_data = 12'h000;
			{8'd166, 8'd68}: color_data = 12'h000;
			{8'd166, 8'd69}: color_data = 12'h000;
			{8'd166, 8'd70}: color_data = 12'h000;
			{8'd166, 8'd71}: color_data = 12'h000;
			{8'd167, 8'd68}: color_data = 12'h000;
			{8'd167, 8'd69}: color_data = 12'h000;
			{8'd167, 8'd70}: color_data = 12'h000;
			{8'd167, 8'd71}: color_data = 12'h000;
			{8'd168, 8'd67}: color_data = 12'h000;
			{8'd168, 8'd68}: color_data = 12'h000;
			{8'd168, 8'd69}: color_data = 12'h000;
			{8'd168, 8'd70}: color_data = 12'h000;
			{8'd168, 8'd71}: color_data = 12'h000;
			{8'd168, 8'd72}: color_data = 12'h000;
			{8'd169, 8'd67}: color_data = 12'h000;
			{8'd169, 8'd68}: color_data = 12'h000;
			{8'd169, 8'd69}: color_data = 12'h000;
			{8'd169, 8'd70}: color_data = 12'h000;
			{8'd169, 8'd71}: color_data = 12'h000;
			{8'd169, 8'd72}: color_data = 12'h000;
            default: color_data = 12'h3b9;
        endcase
endmodule   
