module game_over_rom(
        input wire clk,
        input wire [7:0] x,
        input wire [7:0] y,
        output reg [11:0] color_data
);

    (* rom_style = "block" *)

    //signal declaration
    reg [7:0] x_reg;
    reg [7:0] y_reg;

    always @(posedge clk) begin
        x_reg <= x;
        y_reg <= y;
    end

    always @*
        case ({x_reg, y_reg})
			// right: 8'd235, bottom: 8'd159
			{8'd12, 8'd39}: color_data = 12'h931;
			{8'd12, 8'd40}: color_data = 12'h930;
			{8'd12, 8'd41}: color_data = 12'h930;
			{8'd12, 8'd42}: color_data = 12'h830;
			{8'd12, 8'd43}: color_data = 12'h830;
			{8'd12, 8'd44}: color_data = 12'h830;
			{8'd12, 8'd45}: color_data = 12'h840;
			{8'd12, 8'd46}: color_data = 12'h740;
			{8'd12, 8'd47}: color_data = 12'h700;
			{8'd13, 8'd37}: color_data = 12'h000;
			{8'd13, 8'd38}: color_data = 12'ha30;
			{8'd13, 8'd39}: color_data = 12'hb31;
			{8'd13, 8'd40}: color_data = 12'hb41;
			{8'd13, 8'd41}: color_data = 12'hb41;
			{8'd13, 8'd42}: color_data = 12'hb41;
			{8'd13, 8'd43}: color_data = 12'ha40;
			{8'd13, 8'd44}: color_data = 12'ha50;
			{8'd13, 8'd45}: color_data = 12'ha50;
			{8'd13, 8'd46}: color_data = 12'ha50;
			{8'd13, 8'd47}: color_data = 12'ha50;
			{8'd13, 8'd48}: color_data = 12'ha50;
			{8'd14, 8'd36}: color_data = 12'h300;
			{8'd14, 8'd37}: color_data = 12'ha31;
			{8'd14, 8'd38}: color_data = 12'hc31;
			{8'd14, 8'd39}: color_data = 12'he41;
			{8'd14, 8'd40}: color_data = 12'he51;
			{8'd14, 8'd41}: color_data = 12'he51;
			{8'd14, 8'd42}: color_data = 12'hd61;
			{8'd14, 8'd43}: color_data = 12'hd61;
			{8'd14, 8'd44}: color_data = 12'hd61;
			{8'd14, 8'd45}: color_data = 12'hd71;
			{8'd14, 8'd46}: color_data = 12'hd71;
			{8'd14, 8'd47}: color_data = 12'hd70;
			{8'd14, 8'd48}: color_data = 12'hc60;
			{8'd14, 8'd49}: color_data = 12'ha60;
			{8'd15, 8'd35}: color_data = 12'h000;
			{8'd15, 8'd36}: color_data = 12'hb21;
			{8'd15, 8'd37}: color_data = 12'hc31;
			{8'd15, 8'd38}: color_data = 12'he41;
			{8'd15, 8'd39}: color_data = 12'he41;
			{8'd15, 8'd40}: color_data = 12'he51;
			{8'd15, 8'd41}: color_data = 12'he51;
			{8'd15, 8'd42}: color_data = 12'he61;
			{8'd15, 8'd43}: color_data = 12'he61;
			{8'd15, 8'd44}: color_data = 12'he71;
			{8'd15, 8'd45}: color_data = 12'he71;
			{8'd15, 8'd46}: color_data = 12'he71;
			{8'd15, 8'd47}: color_data = 12'he80;
			{8'd15, 8'd48}: color_data = 12'hd70;
			{8'd15, 8'd49}: color_data = 12'hb60;
			{8'd15, 8'd50}: color_data = 12'h950;
			{8'd16, 8'd34}: color_data = 12'h910;
			{8'd16, 8'd35}: color_data = 12'ha21;
			{8'd16, 8'd36}: color_data = 12'hd31;
			{8'd16, 8'd37}: color_data = 12'he31;
			{8'd16, 8'd38}: color_data = 12'he41;
			{8'd16, 8'd39}: color_data = 12'he41;
			{8'd16, 8'd40}: color_data = 12'he51;
			{8'd16, 8'd41}: color_data = 12'he51;
			{8'd16, 8'd42}: color_data = 12'he61;
			{8'd16, 8'd43}: color_data = 12'he61;
			{8'd16, 8'd44}: color_data = 12'he61;
			{8'd16, 8'd45}: color_data = 12'he71;
			{8'd16, 8'd46}: color_data = 12'he71;
			{8'd16, 8'd47}: color_data = 12'he70;
			{8'd16, 8'd48}: color_data = 12'he80;
			{8'd16, 8'd49}: color_data = 12'hd80;
			{8'd16, 8'd50}: color_data = 12'hb60;
			{8'd16, 8'd51}: color_data = 12'h850;
			{8'd17, 8'd33}: color_data = 12'h811;
			{8'd17, 8'd34}: color_data = 12'ha11;
			{8'd17, 8'd35}: color_data = 12'hd21;
			{8'd17, 8'd36}: color_data = 12'hd31;
			{8'd17, 8'd37}: color_data = 12'hd31;
			{8'd17, 8'd38}: color_data = 12'he41;
			{8'd17, 8'd39}: color_data = 12'he41;
			{8'd17, 8'd40}: color_data = 12'he51;
			{8'd17, 8'd41}: color_data = 12'he51;
			{8'd17, 8'd42}: color_data = 12'he61;
			{8'd17, 8'd43}: color_data = 12'he61;
			{8'd17, 8'd44}: color_data = 12'he71;
			{8'd17, 8'd45}: color_data = 12'he71;
			{8'd17, 8'd46}: color_data = 12'he71;
			{8'd17, 8'd47}: color_data = 12'he80;
			{8'd17, 8'd48}: color_data = 12'he80;
			{8'd17, 8'd49}: color_data = 12'he80;
			{8'd17, 8'd50}: color_data = 12'hd80;
			{8'd17, 8'd51}: color_data = 12'ha60;
			{8'd17, 8'd52}: color_data = 12'h740;
			{8'd18, 8'd32}: color_data = 12'h801;
			{8'd18, 8'd33}: color_data = 12'hb11;
			{8'd18, 8'd34}: color_data = 12'hd11;
			{8'd18, 8'd35}: color_data = 12'hd21;
			{8'd18, 8'd36}: color_data = 12'hd31;
			{8'd18, 8'd37}: color_data = 12'hd31;
			{8'd18, 8'd38}: color_data = 12'he41;
			{8'd18, 8'd39}: color_data = 12'hc41;
			{8'd18, 8'd40}: color_data = 12'hb40;
			{8'd18, 8'd41}: color_data = 12'hc51;
			{8'd18, 8'd42}: color_data = 12'hd51;
			{8'd18, 8'd43}: color_data = 12'hd61;
			{8'd18, 8'd44}: color_data = 12'hd61;
			{8'd18, 8'd45}: color_data = 12'hd71;
			{8'd18, 8'd46}: color_data = 12'he71;
			{8'd18, 8'd47}: color_data = 12'he80;
			{8'd18, 8'd48}: color_data = 12'he80;
			{8'd18, 8'd49}: color_data = 12'he80;
			{8'd18, 8'd50}: color_data = 12'he90;
			{8'd18, 8'd51}: color_data = 12'hd80;
			{8'd18, 8'd52}: color_data = 12'hb70;
			{8'd18, 8'd53}: color_data = 12'h500;
			{8'd19, 8'd31}: color_data = 12'h801;
			{8'd19, 8'd32}: color_data = 12'ha01;
			{8'd19, 8'd33}: color_data = 12'hd11;
			{8'd19, 8'd34}: color_data = 12'hd11;
			{8'd19, 8'd35}: color_data = 12'hd21;
			{8'd19, 8'd36}: color_data = 12'hd31;
			{8'd19, 8'd37}: color_data = 12'hd31;
			{8'd19, 8'd38}: color_data = 12'hb31;
			{8'd19, 8'd39}: color_data = 12'h920;
			{8'd19, 8'd40}: color_data = 12'h930;
			{8'd19, 8'd41}: color_data = 12'ha30;
			{8'd19, 8'd42}: color_data = 12'hc51;
			{8'd19, 8'd43}: color_data = 12'hd51;
			{8'd19, 8'd44}: color_data = 12'hc61;
			{8'd19, 8'd45}: color_data = 12'hb60;
			{8'd19, 8'd46}: color_data = 12'hd71;
			{8'd19, 8'd47}: color_data = 12'he80;
			{8'd19, 8'd48}: color_data = 12'he80;
			{8'd19, 8'd49}: color_data = 12'he80;
			{8'd19, 8'd50}: color_data = 12'he80;
			{8'd19, 8'd51}: color_data = 12'he90;
			{8'd19, 8'd52}: color_data = 12'hd80;
			{8'd19, 8'd53}: color_data = 12'hb70;
			{8'd20, 8'd30}: color_data = 12'h901;
			{8'd20, 8'd31}: color_data = 12'ha01;
			{8'd20, 8'd32}: color_data = 12'hd01;
			{8'd20, 8'd33}: color_data = 12'hd11;
			{8'd20, 8'd34}: color_data = 12'hd11;
			{8'd20, 8'd35}: color_data = 12'hd21;
			{8'd20, 8'd36}: color_data = 12'hd31;
			{8'd20, 8'd37}: color_data = 12'hc31;
			{8'd20, 8'd38}: color_data = 12'h930;
			{8'd20, 8'd45}: color_data = 12'ha51;
			{8'd20, 8'd46}: color_data = 12'hb50;
			{8'd20, 8'd47}: color_data = 12'hc70;
			{8'd20, 8'd48}: color_data = 12'he80;
			{8'd20, 8'd49}: color_data = 12'he80;
			{8'd20, 8'd50}: color_data = 12'he80;
			{8'd20, 8'd51}: color_data = 12'he90;
			{8'd20, 8'd52}: color_data = 12'he90;
			{8'd20, 8'd53}: color_data = 12'hc80;
			{8'd20, 8'd54}: color_data = 12'hf00;
			{8'd21, 8'd29}: color_data = 12'h701;
			{8'd21, 8'd30}: color_data = 12'hb01;
			{8'd21, 8'd31}: color_data = 12'hd01;
			{8'd21, 8'd32}: color_data = 12'hd01;
			{8'd21, 8'd33}: color_data = 12'hd11;
			{8'd21, 8'd34}: color_data = 12'hd11;
			{8'd21, 8'd35}: color_data = 12'hd21;
			{8'd21, 8'd36}: color_data = 12'hc21;
			{8'd21, 8'd37}: color_data = 12'hb21;
			{8'd21, 8'd47}: color_data = 12'hc60;
			{8'd21, 8'd48}: color_data = 12'hd80;
			{8'd21, 8'd49}: color_data = 12'he80;
			{8'd21, 8'd50}: color_data = 12'he80;
			{8'd21, 8'd51}: color_data = 12'he90;
			{8'd21, 8'd52}: color_data = 12'he90;
			{8'd21, 8'd53}: color_data = 12'hd90;
			{8'd21, 8'd54}: color_data = 12'hff0;
			{8'd22, 8'd29}: color_data = 12'ha01;
			{8'd22, 8'd30}: color_data = 12'hc02;
			{8'd22, 8'd31}: color_data = 12'hd02;
			{8'd22, 8'd32}: color_data = 12'hd01;
			{8'd22, 8'd33}: color_data = 12'hd11;
			{8'd22, 8'd34}: color_data = 12'hd11;
			{8'd22, 8'd35}: color_data = 12'hb21;
			{8'd22, 8'd36}: color_data = 12'ha10;
			{8'd22, 8'd47}: color_data = 12'hd70;
			{8'd22, 8'd48}: color_data = 12'hd80;
			{8'd22, 8'd49}: color_data = 12'he80;
			{8'd22, 8'd50}: color_data = 12'he80;
			{8'd22, 8'd51}: color_data = 12'he90;
			{8'd22, 8'd52}: color_data = 12'he90;
			{8'd22, 8'd53}: color_data = 12'hd90;
			{8'd22, 8'd54}: color_data = 12'hff0;
			{8'd23, 8'd29}: color_data = 12'ha01;
			{8'd23, 8'd30}: color_data = 12'hc02;
			{8'd23, 8'd31}: color_data = 12'hd02;
			{8'd23, 8'd32}: color_data = 12'hd01;
			{8'd23, 8'd33}: color_data = 12'hd11;
			{8'd23, 8'd34}: color_data = 12'hb11;
			{8'd23, 8'd35}: color_data = 12'h910;
			{8'd23, 8'd40}: color_data = 12'h000;
			{8'd23, 8'd41}: color_data = 12'h000;
			{8'd23, 8'd42}: color_data = 12'h000;
			{8'd23, 8'd47}: color_data = 12'hc70;
			{8'd23, 8'd48}: color_data = 12'hd80;
			{8'd23, 8'd49}: color_data = 12'he80;
			{8'd23, 8'd50}: color_data = 12'he80;
			{8'd23, 8'd51}: color_data = 12'he90;
			{8'd23, 8'd52}: color_data = 12'he90;
			{8'd23, 8'd53}: color_data = 12'hd90;
			{8'd23, 8'd54}: color_data = 12'hff0;
			{8'd24, 8'd29}: color_data = 12'hb02;
			{8'd24, 8'd30}: color_data = 12'hc02;
			{8'd24, 8'd31}: color_data = 12'hd01;
			{8'd24, 8'd32}: color_data = 12'hd01;
			{8'd24, 8'd33}: color_data = 12'hd11;
			{8'd24, 8'd34}: color_data = 12'hb11;
			{8'd24, 8'd35}: color_data = 12'h810;
			{8'd24, 8'd38}: color_data = 12'ha50;
			{8'd24, 8'd39}: color_data = 12'h930;
			{8'd24, 8'd40}: color_data = 12'h930;
			{8'd24, 8'd41}: color_data = 12'ha40;
			{8'd24, 8'd42}: color_data = 12'hb40;
			{8'd24, 8'd43}: color_data = 12'ha40;
			{8'd24, 8'd44}: color_data = 12'ha30;
			{8'd24, 8'd47}: color_data = 12'hc70;
			{8'd24, 8'd48}: color_data = 12'hd80;
			{8'd24, 8'd49}: color_data = 12'he80;
			{8'd24, 8'd50}: color_data = 12'he80;
			{8'd24, 8'd51}: color_data = 12'he90;
			{8'd24, 8'd52}: color_data = 12'he90;
			{8'd24, 8'd53}: color_data = 12'hd90;
			{8'd24, 8'd54}: color_data = 12'hff0;
			{8'd25, 8'd29}: color_data = 12'hc02;
			{8'd25, 8'd30}: color_data = 12'hd02;
			{8'd25, 8'd31}: color_data = 12'hd01;
			{8'd25, 8'd32}: color_data = 12'hd01;
			{8'd25, 8'd33}: color_data = 12'hd11;
			{8'd25, 8'd34}: color_data = 12'hc11;
			{8'd25, 8'd35}: color_data = 12'ha11;
			{8'd25, 8'd36}: color_data = 12'h911;
			{8'd25, 8'd38}: color_data = 12'h831;
			{8'd25, 8'd39}: color_data = 12'hb41;
			{8'd25, 8'd40}: color_data = 12'hd51;
			{8'd25, 8'd41}: color_data = 12'hd51;
			{8'd25, 8'd42}: color_data = 12'hd51;
			{8'd25, 8'd43}: color_data = 12'hb50;
			{8'd25, 8'd44}: color_data = 12'h940;
			{8'd25, 8'd47}: color_data = 12'hc70;
			{8'd25, 8'd48}: color_data = 12'hd80;
			{8'd25, 8'd49}: color_data = 12'he80;
			{8'd25, 8'd50}: color_data = 12'he80;
			{8'd25, 8'd51}: color_data = 12'he90;
			{8'd25, 8'd52}: color_data = 12'he90;
			{8'd25, 8'd53}: color_data = 12'hd90;
			{8'd25, 8'd54}: color_data = 12'hff0;
			{8'd26, 8'd29}: color_data = 12'hb02;
			{8'd26, 8'd30}: color_data = 12'hd02;
			{8'd26, 8'd31}: color_data = 12'hd01;
			{8'd26, 8'd32}: color_data = 12'hd01;
			{8'd26, 8'd33}: color_data = 12'hd11;
			{8'd26, 8'd34}: color_data = 12'hd11;
			{8'd26, 8'd35}: color_data = 12'hd21;
			{8'd26, 8'd36}: color_data = 12'hb21;
			{8'd26, 8'd37}: color_data = 12'h933;
			{8'd26, 8'd38}: color_data = 12'h730;
			{8'd26, 8'd39}: color_data = 12'hd41;
			{8'd26, 8'd40}: color_data = 12'he51;
			{8'd26, 8'd41}: color_data = 12'he51;
			{8'd26, 8'd42}: color_data = 12'he61;
			{8'd26, 8'd43}: color_data = 12'hc51;
			{8'd26, 8'd44}: color_data = 12'ha40;
			{8'd26, 8'd47}: color_data = 12'hc70;
			{8'd26, 8'd48}: color_data = 12'hd80;
			{8'd26, 8'd49}: color_data = 12'he80;
			{8'd26, 8'd50}: color_data = 12'he80;
			{8'd26, 8'd51}: color_data = 12'he90;
			{8'd26, 8'd52}: color_data = 12'he90;
			{8'd26, 8'd53}: color_data = 12'he90;
			{8'd26, 8'd54}: color_data = 12'hff0;
			{8'd27, 8'd29}: color_data = 12'ha01;
			{8'd27, 8'd30}: color_data = 12'hb02;
			{8'd27, 8'd31}: color_data = 12'hd01;
			{8'd27, 8'd32}: color_data = 12'hd01;
			{8'd27, 8'd33}: color_data = 12'hd11;
			{8'd27, 8'd34}: color_data = 12'hd11;
			{8'd27, 8'd35}: color_data = 12'hd21;
			{8'd27, 8'd36}: color_data = 12'hc21;
			{8'd27, 8'd39}: color_data = 12'hd41;
			{8'd27, 8'd40}: color_data = 12'he51;
			{8'd27, 8'd41}: color_data = 12'he51;
			{8'd27, 8'd42}: color_data = 12'he61;
			{8'd27, 8'd43}: color_data = 12'hc51;
			{8'd27, 8'd44}: color_data = 12'h940;
			{8'd27, 8'd46}: color_data = 12'h330;
			{8'd27, 8'd47}: color_data = 12'hc60;
			{8'd27, 8'd48}: color_data = 12'hd80;
			{8'd27, 8'd49}: color_data = 12'he80;
			{8'd27, 8'd50}: color_data = 12'he80;
			{8'd27, 8'd51}: color_data = 12'he90;
			{8'd27, 8'd52}: color_data = 12'he90;
			{8'd27, 8'd53}: color_data = 12'hd80;
			{8'd27, 8'd54}: color_data = 12'h000;
			{8'd28, 8'd30}: color_data = 12'ha01;
			{8'd28, 8'd31}: color_data = 12'hb01;
			{8'd28, 8'd32}: color_data = 12'hd01;
			{8'd28, 8'd33}: color_data = 12'hd11;
			{8'd28, 8'd34}: color_data = 12'he11;
			{8'd28, 8'd35}: color_data = 12'he21;
			{8'd28, 8'd36}: color_data = 12'hc21;
			{8'd28, 8'd38}: color_data = 12'h200;
			{8'd28, 8'd39}: color_data = 12'hc41;
			{8'd28, 8'd40}: color_data = 12'he51;
			{8'd28, 8'd41}: color_data = 12'he51;
			{8'd28, 8'd42}: color_data = 12'he61;
			{8'd28, 8'd43}: color_data = 12'hc51;
			{8'd28, 8'd44}: color_data = 12'h940;
			{8'd28, 8'd45}: color_data = 12'ha51;
			{8'd28, 8'd46}: color_data = 12'hb60;
			{8'd28, 8'd47}: color_data = 12'hd70;
			{8'd28, 8'd48}: color_data = 12'he80;
			{8'd28, 8'd49}: color_data = 12'he80;
			{8'd28, 8'd50}: color_data = 12'he90;
			{8'd28, 8'd51}: color_data = 12'he90;
			{8'd28, 8'd52}: color_data = 12'hc80;
			{8'd28, 8'd53}: color_data = 12'ha60;
			{8'd29, 8'd31}: color_data = 12'h901;
			{8'd29, 8'd32}: color_data = 12'ha01;
			{8'd29, 8'd33}: color_data = 12'hb11;
			{8'd29, 8'd34}: color_data = 12'hb11;
			{8'd29, 8'd35}: color_data = 12'hb21;
			{8'd29, 8'd36}: color_data = 12'hd31;
			{8'd29, 8'd38}: color_data = 12'h620;
			{8'd29, 8'd39}: color_data = 12'hb40;
			{8'd29, 8'd40}: color_data = 12'he51;
			{8'd29, 8'd41}: color_data = 12'he51;
			{8'd29, 8'd42}: color_data = 12'he61;
			{8'd29, 8'd43}: color_data = 12'he61;
			{8'd29, 8'd44}: color_data = 12'hd61;
			{8'd29, 8'd45}: color_data = 12'hd61;
			{8'd29, 8'd46}: color_data = 12'he71;
			{8'd29, 8'd47}: color_data = 12'he80;
			{8'd29, 8'd48}: color_data = 12'he80;
			{8'd29, 8'd49}: color_data = 12'he80;
			{8'd29, 8'd50}: color_data = 12'he90;
			{8'd29, 8'd51}: color_data = 12'hc80;
			{8'd29, 8'd52}: color_data = 12'h850;
			{8'd29, 8'd53}: color_data = 12'h530;
			{8'd30, 8'd32}: color_data = 12'h900;
			{8'd30, 8'd33}: color_data = 12'h910;
			{8'd30, 8'd34}: color_data = 12'h800;
			{8'd30, 8'd35}: color_data = 12'h810;
			{8'd30, 8'd38}: color_data = 12'h720;
			{8'd30, 8'd39}: color_data = 12'hc41;
			{8'd30, 8'd40}: color_data = 12'he51;
			{8'd30, 8'd41}: color_data = 12'he51;
			{8'd30, 8'd42}: color_data = 12'he61;
			{8'd30, 8'd43}: color_data = 12'he61;
			{8'd30, 8'd44}: color_data = 12'he71;
			{8'd30, 8'd45}: color_data = 12'he71;
			{8'd30, 8'd46}: color_data = 12'he71;
			{8'd30, 8'd47}: color_data = 12'he80;
			{8'd30, 8'd48}: color_data = 12'he80;
			{8'd30, 8'd49}: color_data = 12'he80;
			{8'd30, 8'd50}: color_data = 12'hc70;
			{8'd30, 8'd51}: color_data = 12'h960;
			{8'd30, 8'd52}: color_data = 12'h000;
			{8'd31, 8'd38}: color_data = 12'ha20;
			{8'd31, 8'd39}: color_data = 12'hb40;
			{8'd31, 8'd40}: color_data = 12'hc41;
			{8'd31, 8'd41}: color_data = 12'hc41;
			{8'd31, 8'd42}: color_data = 12'hb41;
			{8'd31, 8'd43}: color_data = 12'hb51;
			{8'd31, 8'd44}: color_data = 12'hb50;
			{8'd31, 8'd45}: color_data = 12'hc61;
			{8'd31, 8'd46}: color_data = 12'hd71;
			{8'd31, 8'd47}: color_data = 12'hd70;
			{8'd31, 8'd48}: color_data = 12'hd70;
			{8'd31, 8'd49}: color_data = 12'hb70;
			{8'd31, 8'd50}: color_data = 12'ha60;
			{8'd32, 8'd39}: color_data = 12'ha30;
			{8'd32, 8'd40}: color_data = 12'ha30;
			{8'd32, 8'd41}: color_data = 12'h930;
			{8'd32, 8'd42}: color_data = 12'h940;
			{8'd32, 8'd43}: color_data = 12'h940;
			{8'd32, 8'd44}: color_data = 12'h930;
			{8'd32, 8'd45}: color_data = 12'h840;
			{8'd32, 8'd46}: color_data = 12'hb60;
			{8'd32, 8'd47}: color_data = 12'hb60;
			{8'd32, 8'd48}: color_data = 12'h960;
			{8'd32, 8'd49}: color_data = 12'h850;
			{8'd32, 8'd50}: color_data = 12'h000;
			{8'd37, 8'd49}: color_data = 12'h940;
			{8'd37, 8'd50}: color_data = 12'hb70;
			{8'd37, 8'd51}: color_data = 12'hc80;
			{8'd37, 8'd52}: color_data = 12'hc80;
			{8'd38, 8'd46}: color_data = 12'h000;
			{8'd38, 8'd47}: color_data = 12'h950;
			{8'd38, 8'd48}: color_data = 12'ha60;
			{8'd38, 8'd49}: color_data = 12'hc70;
			{8'd38, 8'd50}: color_data = 12'hd80;
			{8'd38, 8'd51}: color_data = 12'hd90;
			{8'd38, 8'd52}: color_data = 12'hd80;
			{8'd39, 8'd46}: color_data = 12'ha50;
			{8'd39, 8'd47}: color_data = 12'hb70;
			{8'd39, 8'd48}: color_data = 12'hd80;
			{8'd39, 8'd49}: color_data = 12'he90;
			{8'd39, 8'd50}: color_data = 12'he90;
			{8'd39, 8'd51}: color_data = 12'hd90;
			{8'd39, 8'd52}: color_data = 12'hd90;
			{8'd40, 8'd43}: color_data = 12'h750;
			{8'd40, 8'd44}: color_data = 12'ha50;
			{8'd40, 8'd45}: color_data = 12'hb60;
			{8'd40, 8'd46}: color_data = 12'hc70;
			{8'd40, 8'd47}: color_data = 12'he80;
			{8'd40, 8'd48}: color_data = 12'he80;
			{8'd40, 8'd49}: color_data = 12'he90;
			{8'd40, 8'd50}: color_data = 12'he90;
			{8'd40, 8'd51}: color_data = 12'hd90;
			{8'd40, 8'd52}: color_data = 12'hd90;
			{8'd41, 8'd41}: color_data = 12'ha51;
			{8'd41, 8'd42}: color_data = 12'ha50;
			{8'd41, 8'd43}: color_data = 12'hb50;
			{8'd41, 8'd44}: color_data = 12'hc61;
			{8'd41, 8'd45}: color_data = 12'hd71;
			{8'd41, 8'd46}: color_data = 12'he80;
			{8'd41, 8'd47}: color_data = 12'he80;
			{8'd41, 8'd48}: color_data = 12'he80;
			{8'd41, 8'd49}: color_data = 12'he90;
			{8'd41, 8'd50}: color_data = 12'he90;
			{8'd41, 8'd51}: color_data = 12'hd90;
			{8'd41, 8'd52}: color_data = 12'hd90;
			{8'd42, 8'd39}: color_data = 12'h000;
			{8'd42, 8'd40}: color_data = 12'ha40;
			{8'd42, 8'd41}: color_data = 12'hb41;
			{8'd42, 8'd42}: color_data = 12'hc51;
			{8'd42, 8'd43}: color_data = 12'hd61;
			{8'd42, 8'd44}: color_data = 12'he71;
			{8'd42, 8'd45}: color_data = 12'he71;
			{8'd42, 8'd46}: color_data = 12'he80;
			{8'd42, 8'd47}: color_data = 12'he80;
			{8'd42, 8'd48}: color_data = 12'he80;
			{8'd42, 8'd49}: color_data = 12'he90;
			{8'd42, 8'd50}: color_data = 12'he90;
			{8'd42, 8'd51}: color_data = 12'hd90;
			{8'd42, 8'd52}: color_data = 12'hd90;
			{8'd43, 8'd37}: color_data = 12'h502;
			{8'd43, 8'd38}: color_data = 12'ha30;
			{8'd43, 8'd39}: color_data = 12'hb41;
			{8'd43, 8'd40}: color_data = 12'hc51;
			{8'd43, 8'd41}: color_data = 12'he61;
			{8'd43, 8'd42}: color_data = 12'he61;
			{8'd43, 8'd43}: color_data = 12'he71;
			{8'd43, 8'd44}: color_data = 12'he71;
			{8'd43, 8'd45}: color_data = 12'he71;
			{8'd43, 8'd46}: color_data = 12'he80;
			{8'd43, 8'd47}: color_data = 12'he80;
			{8'd43, 8'd48}: color_data = 12'he80;
			{8'd43, 8'd49}: color_data = 12'he90;
			{8'd43, 8'd50}: color_data = 12'he90;
			{8'd43, 8'd51}: color_data = 12'hd90;
			{8'd43, 8'd52}: color_data = 12'hd90;
			{8'd44, 8'd36}: color_data = 12'h930;
			{8'd44, 8'd37}: color_data = 12'hb31;
			{8'd44, 8'd38}: color_data = 12'hc41;
			{8'd44, 8'd39}: color_data = 12'hd51;
			{8'd44, 8'd40}: color_data = 12'he51;
			{8'd44, 8'd41}: color_data = 12'he61;
			{8'd44, 8'd42}: color_data = 12'he61;
			{8'd44, 8'd43}: color_data = 12'he71;
			{8'd44, 8'd44}: color_data = 12'he71;
			{8'd44, 8'd45}: color_data = 12'he71;
			{8'd44, 8'd46}: color_data = 12'he80;
			{8'd44, 8'd47}: color_data = 12'he80;
			{8'd44, 8'd48}: color_data = 12'he80;
			{8'd44, 8'd49}: color_data = 12'he90;
			{8'd44, 8'd50}: color_data = 12'he90;
			{8'd44, 8'd51}: color_data = 12'hd90;
			{8'd44, 8'd52}: color_data = 12'hc80;
			{8'd45, 8'd33}: color_data = 12'hf00;
			{8'd45, 8'd34}: color_data = 12'h921;
			{8'd45, 8'd35}: color_data = 12'hb20;
			{8'd45, 8'd36}: color_data = 12'hc31;
			{8'd45, 8'd37}: color_data = 12'hd41;
			{8'd45, 8'd38}: color_data = 12'he41;
			{8'd45, 8'd39}: color_data = 12'he51;
			{8'd45, 8'd40}: color_data = 12'he51;
			{8'd45, 8'd41}: color_data = 12'he61;
			{8'd45, 8'd42}: color_data = 12'he61;
			{8'd45, 8'd43}: color_data = 12'he71;
			{8'd45, 8'd44}: color_data = 12'he71;
			{8'd45, 8'd45}: color_data = 12'he71;
			{8'd45, 8'd46}: color_data = 12'he80;
			{8'd45, 8'd47}: color_data = 12'he80;
			{8'd45, 8'd48}: color_data = 12'hd80;
			{8'd45, 8'd49}: color_data = 12'hc80;
			{8'd45, 8'd50}: color_data = 12'hd90;
			{8'd45, 8'd51}: color_data = 12'hc80;
			{8'd45, 8'd52}: color_data = 12'h960;
			{8'd46, 8'd31}: color_data = 12'hf00;
			{8'd46, 8'd32}: color_data = 12'ha01;
			{8'd46, 8'd33}: color_data = 12'hb11;
			{8'd46, 8'd34}: color_data = 12'hc11;
			{8'd46, 8'd35}: color_data = 12'hd21;
			{8'd46, 8'd36}: color_data = 12'he31;
			{8'd46, 8'd37}: color_data = 12'he41;
			{8'd46, 8'd38}: color_data = 12'he41;
			{8'd46, 8'd39}: color_data = 12'he51;
			{8'd46, 8'd40}: color_data = 12'he51;
			{8'd46, 8'd41}: color_data = 12'hd51;
			{8'd46, 8'd42}: color_data = 12'hb50;
			{8'd46, 8'd43}: color_data = 12'hb50;
			{8'd46, 8'd44}: color_data = 12'hd61;
			{8'd46, 8'd45}: color_data = 12'he71;
			{8'd46, 8'd46}: color_data = 12'he80;
			{8'd46, 8'd47}: color_data = 12'hd70;
			{8'd46, 8'd48}: color_data = 12'ha60;
			{8'd46, 8'd49}: color_data = 12'ha60;
			{8'd46, 8'd50}: color_data = 12'ha70;
			{8'd46, 8'd51}: color_data = 12'ha70;
			{8'd46, 8'd52}: color_data = 12'h971;
			{8'd47, 8'd31}: color_data = 12'ha01;
			{8'd47, 8'd32}: color_data = 12'hb01;
			{8'd47, 8'd33}: color_data = 12'hd11;
			{8'd47, 8'd34}: color_data = 12'hd21;
			{8'd47, 8'd35}: color_data = 12'hd31;
			{8'd47, 8'd36}: color_data = 12'hd31;
			{8'd47, 8'd37}: color_data = 12'hd41;
			{8'd47, 8'd38}: color_data = 12'hd41;
			{8'd47, 8'd39}: color_data = 12'hc41;
			{8'd47, 8'd40}: color_data = 12'hb40;
			{8'd47, 8'd41}: color_data = 12'ha40;
			{8'd47, 8'd42}: color_data = 12'ha40;
			{8'd47, 8'd43}: color_data = 12'h520;
			{8'd47, 8'd44}: color_data = 12'hc61;
			{8'd47, 8'd45}: color_data = 12'he71;
			{8'd47, 8'd46}: color_data = 12'he80;
			{8'd47, 8'd47}: color_data = 12'hc70;
			{8'd47, 8'd48}: color_data = 12'ha60;
			{8'd47, 8'd49}: color_data = 12'h00f;
			{8'd47, 8'd50}: color_data = 12'ha70;
			{8'd47, 8'd51}: color_data = 12'hf00;
			{8'd48, 8'd30}: color_data = 12'h900;
			{8'd48, 8'd31}: color_data = 12'hc01;
			{8'd48, 8'd32}: color_data = 12'hd01;
			{8'd48, 8'd33}: color_data = 12'hd11;
			{8'd48, 8'd34}: color_data = 12'hd21;
			{8'd48, 8'd35}: color_data = 12'hd31;
			{8'd48, 8'd36}: color_data = 12'hd31;
			{8'd48, 8'd37}: color_data = 12'hc31;
			{8'd48, 8'd38}: color_data = 12'ha31;
			{8'd48, 8'd39}: color_data = 12'ha31;
			{8'd48, 8'd40}: color_data = 12'h930;
			{8'd48, 8'd44}: color_data = 12'hd71;
			{8'd48, 8'd45}: color_data = 12'he71;
			{8'd48, 8'd46}: color_data = 12'he80;
			{8'd48, 8'd47}: color_data = 12'hd80;
			{8'd48, 8'd48}: color_data = 12'hc70;
			{8'd49, 8'd30}: color_data = 12'hb01;
			{8'd49, 8'd31}: color_data = 12'hc01;
			{8'd49, 8'd32}: color_data = 12'hd01;
			{8'd49, 8'd33}: color_data = 12'hd11;
			{8'd49, 8'd34}: color_data = 12'hd21;
			{8'd49, 8'd35}: color_data = 12'hd31;
			{8'd49, 8'd36}: color_data = 12'hd31;
			{8'd49, 8'd37}: color_data = 12'hb31;
			{8'd49, 8'd38}: color_data = 12'h820;
			{8'd49, 8'd44}: color_data = 12'hd71;
			{8'd49, 8'd45}: color_data = 12'he71;
			{8'd49, 8'd46}: color_data = 12'he80;
			{8'd49, 8'd47}: color_data = 12'he80;
			{8'd49, 8'd48}: color_data = 12'hc70;
			{8'd49, 8'd49}: color_data = 12'h930;
			{8'd50, 8'd31}: color_data = 12'hb01;
			{8'd50, 8'd32}: color_data = 12'hd01;
			{8'd50, 8'd33}: color_data = 12'hd11;
			{8'd50, 8'd34}: color_data = 12'hd21;
			{8'd50, 8'd35}: color_data = 12'hd31;
			{8'd50, 8'd36}: color_data = 12'hd31;
			{8'd50, 8'd37}: color_data = 12'hc31;
			{8'd50, 8'd38}: color_data = 12'h920;
			{8'd50, 8'd39}: color_data = 12'h622;
			{8'd50, 8'd44}: color_data = 12'hd71;
			{8'd50, 8'd45}: color_data = 12'hd71;
			{8'd50, 8'd46}: color_data = 12'he80;
			{8'd50, 8'd47}: color_data = 12'he80;
			{8'd50, 8'd48}: color_data = 12'hd80;
			{8'd50, 8'd49}: color_data = 12'ha60;
			{8'd50, 8'd50}: color_data = 12'hb70;
			{8'd50, 8'd51}: color_data = 12'hd91;
			{8'd51, 8'd31}: color_data = 12'ha01;
			{8'd51, 8'd32}: color_data = 12'hc01;
			{8'd51, 8'd33}: color_data = 12'hd11;
			{8'd51, 8'd34}: color_data = 12'hd21;
			{8'd51, 8'd35}: color_data = 12'hd31;
			{8'd51, 8'd36}: color_data = 12'hd31;
			{8'd51, 8'd37}: color_data = 12'he41;
			{8'd51, 8'd38}: color_data = 12'hc41;
			{8'd51, 8'd39}: color_data = 12'ha30;
			{8'd51, 8'd40}: color_data = 12'hc41;
			{8'd51, 8'd41}: color_data = 12'hd51;
			{8'd51, 8'd42}: color_data = 12'hd61;
			{8'd51, 8'd43}: color_data = 12'he61;
			{8'd51, 8'd44}: color_data = 12'hd71;
			{8'd51, 8'd45}: color_data = 12'he81;
			{8'd51, 8'd46}: color_data = 12'he80;
			{8'd51, 8'd47}: color_data = 12'he80;
			{8'd51, 8'd48}: color_data = 12'he80;
			{8'd51, 8'd49}: color_data = 12'hd80;
			{8'd51, 8'd50}: color_data = 12'hd90;
			{8'd51, 8'd51}: color_data = 12'he90;
			{8'd51, 8'd52}: color_data = 12'hd80;
			{8'd52, 8'd31}: color_data = 12'h801;
			{8'd52, 8'd32}: color_data = 12'ha01;
			{8'd52, 8'd33}: color_data = 12'hc11;
			{8'd52, 8'd34}: color_data = 12'hd21;
			{8'd52, 8'd35}: color_data = 12'hd31;
			{8'd52, 8'd36}: color_data = 12'hd31;
			{8'd52, 8'd37}: color_data = 12'hd41;
			{8'd52, 8'd38}: color_data = 12'he41;
			{8'd52, 8'd39}: color_data = 12'hd51;
			{8'd52, 8'd40}: color_data = 12'he51;
			{8'd52, 8'd41}: color_data = 12'he61;
			{8'd52, 8'd42}: color_data = 12'he61;
			{8'd52, 8'd43}: color_data = 12'he61;
			{8'd52, 8'd44}: color_data = 12'he71;
			{8'd52, 8'd45}: color_data = 12'he71;
			{8'd52, 8'd46}: color_data = 12'he80;
			{8'd52, 8'd47}: color_data = 12'he80;
			{8'd52, 8'd48}: color_data = 12'he80;
			{8'd52, 8'd49}: color_data = 12'he90;
			{8'd52, 8'd50}: color_data = 12'he90;
			{8'd52, 8'd51}: color_data = 12'he90;
			{8'd52, 8'd52}: color_data = 12'hd90;
			{8'd53, 8'd32}: color_data = 12'h700;
			{8'd53, 8'd33}: color_data = 12'ha11;
			{8'd53, 8'd34}: color_data = 12'hc21;
			{8'd53, 8'd35}: color_data = 12'he31;
			{8'd53, 8'd36}: color_data = 12'hd31;
			{8'd53, 8'd37}: color_data = 12'hd41;
			{8'd53, 8'd38}: color_data = 12'he41;
			{8'd53, 8'd39}: color_data = 12'he51;
			{8'd53, 8'd40}: color_data = 12'he51;
			{8'd53, 8'd41}: color_data = 12'he61;
			{8'd53, 8'd42}: color_data = 12'he61;
			{8'd53, 8'd43}: color_data = 12'he71;
			{8'd53, 8'd44}: color_data = 12'he71;
			{8'd53, 8'd45}: color_data = 12'he71;
			{8'd53, 8'd46}: color_data = 12'he80;
			{8'd53, 8'd47}: color_data = 12'he80;
			{8'd53, 8'd48}: color_data = 12'he80;
			{8'd53, 8'd49}: color_data = 12'he90;
			{8'd53, 8'd50}: color_data = 12'he90;
			{8'd53, 8'd51}: color_data = 12'hd90;
			{8'd53, 8'd52}: color_data = 12'hd90;
			{8'd54, 8'd34}: color_data = 12'ha21;
			{8'd54, 8'd35}: color_data = 12'hc21;
			{8'd54, 8'd36}: color_data = 12'hd31;
			{8'd54, 8'd37}: color_data = 12'he41;
			{8'd54, 8'd38}: color_data = 12'he41;
			{8'd54, 8'd39}: color_data = 12'he51;
			{8'd54, 8'd40}: color_data = 12'he51;
			{8'd54, 8'd41}: color_data = 12'he61;
			{8'd54, 8'd42}: color_data = 12'he61;
			{8'd54, 8'd43}: color_data = 12'he71;
			{8'd54, 8'd44}: color_data = 12'he71;
			{8'd54, 8'd45}: color_data = 12'he71;
			{8'd54, 8'd46}: color_data = 12'he80;
			{8'd54, 8'd47}: color_data = 12'he80;
			{8'd54, 8'd48}: color_data = 12'he80;
			{8'd54, 8'd49}: color_data = 12'he90;
			{8'd54, 8'd50}: color_data = 12'he90;
			{8'd54, 8'd51}: color_data = 12'hd90;
			{8'd54, 8'd52}: color_data = 12'hd90;
			{8'd55, 8'd35}: color_data = 12'ha20;
			{8'd55, 8'd36}: color_data = 12'hc31;
			{8'd55, 8'd37}: color_data = 12'he41;
			{8'd55, 8'd38}: color_data = 12'he41;
			{8'd55, 8'd39}: color_data = 12'he51;
			{8'd55, 8'd40}: color_data = 12'he51;
			{8'd55, 8'd41}: color_data = 12'he61;
			{8'd55, 8'd42}: color_data = 12'he61;
			{8'd55, 8'd43}: color_data = 12'he71;
			{8'd55, 8'd44}: color_data = 12'he71;
			{8'd55, 8'd45}: color_data = 12'he71;
			{8'd55, 8'd46}: color_data = 12'he80;
			{8'd55, 8'd47}: color_data = 12'he80;
			{8'd55, 8'd48}: color_data = 12'he80;
			{8'd55, 8'd49}: color_data = 12'he90;
			{8'd55, 8'd50}: color_data = 12'he90;
			{8'd55, 8'd51}: color_data = 12'hd90;
			{8'd55, 8'd52}: color_data = 12'hd80;
			{8'd56, 8'd36}: color_data = 12'h920;
			{8'd56, 8'd37}: color_data = 12'hb31;
			{8'd56, 8'd38}: color_data = 12'hd41;
			{8'd56, 8'd39}: color_data = 12'he51;
			{8'd56, 8'd40}: color_data = 12'he51;
			{8'd56, 8'd41}: color_data = 12'he61;
			{8'd56, 8'd42}: color_data = 12'he61;
			{8'd56, 8'd43}: color_data = 12'he71;
			{8'd56, 8'd44}: color_data = 12'he71;
			{8'd56, 8'd45}: color_data = 12'he71;
			{8'd56, 8'd46}: color_data = 12'he80;
			{8'd56, 8'd47}: color_data = 12'he80;
			{8'd56, 8'd48}: color_data = 12'he80;
			{8'd56, 8'd49}: color_data = 12'he90;
			{8'd56, 8'd50}: color_data = 12'he90;
			{8'd56, 8'd51}: color_data = 12'hd90;
			{8'd56, 8'd52}: color_data = 12'ha70;
			{8'd57, 8'd37}: color_data = 12'h920;
			{8'd57, 8'd38}: color_data = 12'ha31;
			{8'd57, 8'd39}: color_data = 12'ha31;
			{8'd57, 8'd40}: color_data = 12'ha40;
			{8'd57, 8'd41}: color_data = 12'ha40;
			{8'd57, 8'd42}: color_data = 12'ha50;
			{8'd57, 8'd43}: color_data = 12'ha50;
			{8'd57, 8'd44}: color_data = 12'hb50;
			{8'd57, 8'd45}: color_data = 12'hb60;
			{8'd57, 8'd46}: color_data = 12'hb60;
			{8'd57, 8'd47}: color_data = 12'hb60;
			{8'd57, 8'd48}: color_data = 12'hb70;
			{8'd57, 8'd49}: color_data = 12'hb70;
			{8'd57, 8'd50}: color_data = 12'hb70;
			{8'd57, 8'd51}: color_data = 12'hb70;
			{8'd57, 8'd52}: color_data = 12'h970;
			{8'd58, 8'd38}: color_data = 12'h620;
			{8'd58, 8'd39}: color_data = 12'h820;
			{8'd58, 8'd40}: color_data = 12'h830;
			{8'd58, 8'd41}: color_data = 12'h830;
			{8'd58, 8'd42}: color_data = 12'h830;
			{8'd58, 8'd43}: color_data = 12'h840;
			{8'd58, 8'd44}: color_data = 12'h840;
			{8'd58, 8'd45}: color_data = 12'h940;
			{8'd58, 8'd46}: color_data = 12'h950;
			{8'd58, 8'd47}: color_data = 12'h950;
			{8'd58, 8'd48}: color_data = 12'h950;
			{8'd58, 8'd49}: color_data = 12'h960;
			{8'd58, 8'd50}: color_data = 12'h960;
			{8'd58, 8'd51}: color_data = 12'ha60;
			{8'd58, 8'd52}: color_data = 12'h970;
			{8'd64, 8'd50}: color_data = 12'h850;
			{8'd64, 8'd51}: color_data = 12'ha60;
			{8'd64, 8'd52}: color_data = 12'hc70;
			{8'd64, 8'd53}: color_data = 12'hc70;
			{8'd65, 8'd47}: color_data = 12'h730;
			{8'd65, 8'd48}: color_data = 12'ha60;
			{8'd65, 8'd49}: color_data = 12'hb60;
			{8'd65, 8'd50}: color_data = 12'hb70;
			{8'd65, 8'd51}: color_data = 12'hd80;
			{8'd65, 8'd52}: color_data = 12'hd80;
			{8'd65, 8'd53}: color_data = 12'hc80;
			{8'd66, 8'd45}: color_data = 12'h731;
			{8'd66, 8'd46}: color_data = 12'h940;
			{8'd66, 8'd47}: color_data = 12'hb60;
			{8'd66, 8'd48}: color_data = 12'hc70;
			{8'd66, 8'd49}: color_data = 12'hd70;
			{8'd66, 8'd50}: color_data = 12'he80;
			{8'd66, 8'd51}: color_data = 12'he80;
			{8'd66, 8'd52}: color_data = 12'he90;
			{8'd66, 8'd53}: color_data = 12'hc80;
			{8'd66, 8'd54}: color_data = 12'ha70;
			{8'd67, 8'd38}: color_data = 12'h710;
			{8'd67, 8'd39}: color_data = 12'h810;
			{8'd67, 8'd40}: color_data = 12'h920;
			{8'd67, 8'd41}: color_data = 12'ha30;
			{8'd67, 8'd42}: color_data = 12'hc41;
			{8'd67, 8'd43}: color_data = 12'hd51;
			{8'd67, 8'd44}: color_data = 12'hc51;
			{8'd67, 8'd45}: color_data = 12'ha50;
			{8'd67, 8'd46}: color_data = 12'hc61;
			{8'd67, 8'd47}: color_data = 12'hd71;
			{8'd67, 8'd48}: color_data = 12'he81;
			{8'd67, 8'd49}: color_data = 12'he80;
			{8'd67, 8'd50}: color_data = 12'he80;
			{8'd67, 8'd51}: color_data = 12'he80;
			{8'd67, 8'd52}: color_data = 12'he90;
			{8'd67, 8'd53}: color_data = 12'hd80;
			{8'd67, 8'd54}: color_data = 12'hb70;
			{8'd68, 8'd32}: color_data = 12'h900;
			{8'd68, 8'd33}: color_data = 12'hb01;
			{8'd68, 8'd34}: color_data = 12'hb01;
			{8'd68, 8'd35}: color_data = 12'hd11;
			{8'd68, 8'd36}: color_data = 12'hd21;
			{8'd68, 8'd37}: color_data = 12'hc21;
			{8'd68, 8'd38}: color_data = 12'hb21;
			{8'd68, 8'd39}: color_data = 12'ha21;
			{8'd68, 8'd40}: color_data = 12'hb31;
			{8'd68, 8'd41}: color_data = 12'hc41;
			{8'd68, 8'd42}: color_data = 12'hd51;
			{8'd68, 8'd43}: color_data = 12'he51;
			{8'd68, 8'd44}: color_data = 12'hd61;
			{8'd68, 8'd45}: color_data = 12'hd61;
			{8'd68, 8'd46}: color_data = 12'he61;
			{8'd68, 8'd47}: color_data = 12'he71;
			{8'd68, 8'd48}: color_data = 12'he71;
			{8'd68, 8'd49}: color_data = 12'he80;
			{8'd68, 8'd50}: color_data = 12'he80;
			{8'd68, 8'd51}: color_data = 12'he80;
			{8'd68, 8'd52}: color_data = 12'he90;
			{8'd68, 8'd53}: color_data = 12'he90;
			{8'd68, 8'd54}: color_data = 12'hd80;
			{8'd68, 8'd55}: color_data = 12'ha70;
			{8'd69, 8'd32}: color_data = 12'h900;
			{8'd69, 8'd33}: color_data = 12'hb01;
			{8'd69, 8'd34}: color_data = 12'hd01;
			{8'd69, 8'd35}: color_data = 12'hd11;
			{8'd69, 8'd36}: color_data = 12'hd21;
			{8'd69, 8'd37}: color_data = 12'hd21;
			{8'd69, 8'd38}: color_data = 12'hd31;
			{8'd69, 8'd39}: color_data = 12'hd41;
			{8'd69, 8'd40}: color_data = 12'he41;
			{8'd69, 8'd41}: color_data = 12'he51;
			{8'd69, 8'd42}: color_data = 12'he51;
			{8'd69, 8'd43}: color_data = 12'he51;
			{8'd69, 8'd44}: color_data = 12'he61;
			{8'd69, 8'd45}: color_data = 12'he61;
			{8'd69, 8'd46}: color_data = 12'he61;
			{8'd69, 8'd47}: color_data = 12'he71;
			{8'd69, 8'd48}: color_data = 12'he71;
			{8'd69, 8'd49}: color_data = 12'he80;
			{8'd69, 8'd50}: color_data = 12'he80;
			{8'd69, 8'd51}: color_data = 12'he80;
			{8'd69, 8'd52}: color_data = 12'hc80;
			{8'd69, 8'd53}: color_data = 12'hc80;
			{8'd69, 8'd54}: color_data = 12'hd80;
			{8'd69, 8'd55}: color_data = 12'hb70;
			{8'd70, 8'd33}: color_data = 12'h901;
			{8'd70, 8'd34}: color_data = 12'hb01;
			{8'd70, 8'd35}: color_data = 12'hd11;
			{8'd70, 8'd36}: color_data = 12'hd21;
			{8'd70, 8'd37}: color_data = 12'hd21;
			{8'd70, 8'd38}: color_data = 12'hd31;
			{8'd70, 8'd39}: color_data = 12'hd41;
			{8'd70, 8'd40}: color_data = 12'he41;
			{8'd70, 8'd41}: color_data = 12'he51;
			{8'd70, 8'd42}: color_data = 12'he51;
			{8'd70, 8'd43}: color_data = 12'he51;
			{8'd70, 8'd44}: color_data = 12'he61;
			{8'd70, 8'd45}: color_data = 12'he61;
			{8'd70, 8'd46}: color_data = 12'he61;
			{8'd70, 8'd47}: color_data = 12'hd71;
			{8'd70, 8'd48}: color_data = 12'hc60;
			{8'd70, 8'd49}: color_data = 12'hc60;
			{8'd70, 8'd50}: color_data = 12'hd70;
			{8'd70, 8'd51}: color_data = 12'hb70;
			{8'd70, 8'd52}: color_data = 12'ha60;
			{8'd70, 8'd53}: color_data = 12'h850;
			{8'd70, 8'd54}: color_data = 12'h700;
			{8'd71, 8'd34}: color_data = 12'h901;
			{8'd71, 8'd35}: color_data = 12'hc11;
			{8'd71, 8'd36}: color_data = 12'hd21;
			{8'd71, 8'd37}: color_data = 12'hd21;
			{8'd71, 8'd38}: color_data = 12'hd31;
			{8'd71, 8'd39}: color_data = 12'hd41;
			{8'd71, 8'd40}: color_data = 12'he41;
			{8'd71, 8'd41}: color_data = 12'he51;
			{8'd71, 8'd42}: color_data = 12'he51;
			{8'd71, 8'd43}: color_data = 12'he51;
			{8'd71, 8'd44}: color_data = 12'hc51;
			{8'd71, 8'd45}: color_data = 12'hb50;
			{8'd71, 8'd46}: color_data = 12'hc51;
			{8'd71, 8'd47}: color_data = 12'hc60;
			{8'd71, 8'd48}: color_data = 12'ha50;
			{8'd71, 8'd49}: color_data = 12'h840;
			{8'd72, 8'd35}: color_data = 12'ha10;
			{8'd72, 8'd36}: color_data = 12'hc21;
			{8'd72, 8'd37}: color_data = 12'hd21;
			{8'd72, 8'd38}: color_data = 12'hd31;
			{8'd72, 8'd39}: color_data = 12'hd41;
			{8'd72, 8'd40}: color_data = 12'he41;
			{8'd72, 8'd41}: color_data = 12'he51;
			{8'd72, 8'd42}: color_data = 12'he51;
			{8'd72, 8'd43}: color_data = 12'hd51;
			{8'd72, 8'd44}: color_data = 12'hb40;
			{8'd72, 8'd45}: color_data = 12'h620;
			{8'd73, 8'd35}: color_data = 12'h000;
			{8'd73, 8'd36}: color_data = 12'hb21;
			{8'd73, 8'd37}: color_data = 12'hd21;
			{8'd73, 8'd38}: color_data = 12'hd31;
			{8'd73, 8'd39}: color_data = 12'hd41;
			{8'd73, 8'd40}: color_data = 12'he41;
			{8'd73, 8'd41}: color_data = 12'he51;
			{8'd73, 8'd42}: color_data = 12'he51;
			{8'd73, 8'd43}: color_data = 12'hd51;
			{8'd73, 8'd44}: color_data = 12'hb51;
			{8'd73, 8'd45}: color_data = 12'ha50;
			{8'd73, 8'd46}: color_data = 12'ha50;
			{8'd74, 8'd36}: color_data = 12'ha10;
			{8'd74, 8'd37}: color_data = 12'hb21;
			{8'd74, 8'd38}: color_data = 12'hd31;
			{8'd74, 8'd39}: color_data = 12'hd41;
			{8'd74, 8'd40}: color_data = 12'he41;
			{8'd74, 8'd41}: color_data = 12'he51;
			{8'd74, 8'd42}: color_data = 12'he51;
			{8'd74, 8'd43}: color_data = 12'he51;
			{8'd74, 8'd44}: color_data = 12'hd61;
			{8'd74, 8'd45}: color_data = 12'hd61;
			{8'd74, 8'd46}: color_data = 12'hb50;
			{8'd74, 8'd47}: color_data = 12'hb60;
			{8'd74, 8'd48}: color_data = 12'hb61;
			{8'd75, 8'd37}: color_data = 12'h921;
			{8'd75, 8'd38}: color_data = 12'hc31;
			{8'd75, 8'd39}: color_data = 12'he41;
			{8'd75, 8'd40}: color_data = 12'he41;
			{8'd75, 8'd41}: color_data = 12'he51;
			{8'd75, 8'd42}: color_data = 12'he51;
			{8'd75, 8'd43}: color_data = 12'he51;
			{8'd75, 8'd44}: color_data = 12'he61;
			{8'd75, 8'd45}: color_data = 12'he61;
			{8'd75, 8'd46}: color_data = 12'he61;
			{8'd75, 8'd47}: color_data = 12'hd71;
			{8'd75, 8'd48}: color_data = 12'hc61;
			{8'd75, 8'd49}: color_data = 12'hb51;
			{8'd76, 8'd37}: color_data = 12'h000;
			{8'd76, 8'd38}: color_data = 12'hc31;
			{8'd76, 8'd39}: color_data = 12'he41;
			{8'd76, 8'd40}: color_data = 12'he41;
			{8'd76, 8'd41}: color_data = 12'he51;
			{8'd76, 8'd42}: color_data = 12'he51;
			{8'd76, 8'd43}: color_data = 12'he51;
			{8'd76, 8'd44}: color_data = 12'he61;
			{8'd76, 8'd45}: color_data = 12'he61;
			{8'd76, 8'd46}: color_data = 12'he61;
			{8'd76, 8'd47}: color_data = 12'hc61;
			{8'd76, 8'd48}: color_data = 12'hc60;
			{8'd76, 8'd49}: color_data = 12'hb61;
			{8'd77, 8'd36}: color_data = 12'h700;
			{8'd77, 8'd37}: color_data = 12'hb21;
			{8'd77, 8'd38}: color_data = 12'hd31;
			{8'd77, 8'd39}: color_data = 12'hd41;
			{8'd77, 8'd40}: color_data = 12'he41;
			{8'd77, 8'd41}: color_data = 12'he51;
			{8'd77, 8'd42}: color_data = 12'he51;
			{8'd77, 8'd43}: color_data = 12'he51;
			{8'd77, 8'd44}: color_data = 12'he61;
			{8'd77, 8'd45}: color_data = 12'hc51;
			{8'd77, 8'd46}: color_data = 12'hb50;
			{8'd77, 8'd47}: color_data = 12'ha50;
			{8'd77, 8'd48}: color_data = 12'h730;
			{8'd78, 8'd35}: color_data = 12'h500;
			{8'd78, 8'd36}: color_data = 12'hb11;
			{8'd78, 8'd37}: color_data = 12'hc21;
			{8'd78, 8'd38}: color_data = 12'he31;
			{8'd78, 8'd39}: color_data = 12'hd41;
			{8'd78, 8'd40}: color_data = 12'he41;
			{8'd78, 8'd41}: color_data = 12'he51;
			{8'd78, 8'd42}: color_data = 12'he51;
			{8'd78, 8'd43}: color_data = 12'hd51;
			{8'd78, 8'd44}: color_data = 12'hb40;
			{8'd78, 8'd45}: color_data = 12'ha40;
			{8'd78, 8'd46}: color_data = 12'h840;
			{8'd79, 8'd35}: color_data = 12'hb11;
			{8'd79, 8'd36}: color_data = 12'hc21;
			{8'd79, 8'd37}: color_data = 12'hd21;
			{8'd79, 8'd38}: color_data = 12'hd31;
			{8'd79, 8'd39}: color_data = 12'hd41;
			{8'd79, 8'd40}: color_data = 12'he41;
			{8'd79, 8'd41}: color_data = 12'he51;
			{8'd79, 8'd42}: color_data = 12'he51;
			{8'd79, 8'd43}: color_data = 12'hb41;
			{8'd79, 8'd44}: color_data = 12'h730;
			{8'd79, 8'd130}: color_data = 12'h000;
			{8'd79, 8'd131}: color_data = 12'h000;
			{8'd79, 8'd132}: color_data = 12'h000;
			{8'd80, 8'd33}: color_data = 12'h700;
			{8'd80, 8'd34}: color_data = 12'hb01;
			{8'd80, 8'd35}: color_data = 12'hc11;
			{8'd80, 8'd36}: color_data = 12'hd21;
			{8'd80, 8'd37}: color_data = 12'hd21;
			{8'd80, 8'd38}: color_data = 12'hd31;
			{8'd80, 8'd39}: color_data = 12'hd41;
			{8'd80, 8'd40}: color_data = 12'he41;
			{8'd80, 8'd41}: color_data = 12'he51;
			{8'd80, 8'd42}: color_data = 12'he51;
			{8'd80, 8'd43}: color_data = 12'hd51;
			{8'd80, 8'd44}: color_data = 12'hd51;
			{8'd80, 8'd45}: color_data = 12'he61;
			{8'd80, 8'd46}: color_data = 12'he61;
			{8'd80, 8'd47}: color_data = 12'he71;
			{8'd80, 8'd48}: color_data = 12'he71;
			{8'd80, 8'd49}: color_data = 12'he70;
			{8'd80, 8'd50}: color_data = 12'he80;
			{8'd80, 8'd51}: color_data = 12'he80;
			{8'd80, 8'd52}: color_data = 12'hd80;
			{8'd80, 8'd53}: color_data = 12'he80;
			{8'd80, 8'd128}: color_data = 12'h000;
			{8'd80, 8'd129}: color_data = 12'h000;
			{8'd80, 8'd130}: color_data = 12'h000;
			{8'd80, 8'd131}: color_data = 12'h000;
			{8'd80, 8'd132}: color_data = 12'h000;
			{8'd80, 8'd133}: color_data = 12'h333;
			{8'd81, 8'd32}: color_data = 12'h700;
			{8'd81, 8'd33}: color_data = 12'hb01;
			{8'd81, 8'd34}: color_data = 12'hc01;
			{8'd81, 8'd35}: color_data = 12'hd11;
			{8'd81, 8'd36}: color_data = 12'hd21;
			{8'd81, 8'd37}: color_data = 12'hd21;
			{8'd81, 8'd38}: color_data = 12'hd31;
			{8'd81, 8'd39}: color_data = 12'hd41;
			{8'd81, 8'd40}: color_data = 12'he41;
			{8'd81, 8'd41}: color_data = 12'he51;
			{8'd81, 8'd42}: color_data = 12'he51;
			{8'd81, 8'd43}: color_data = 12'he51;
			{8'd81, 8'd44}: color_data = 12'he61;
			{8'd81, 8'd45}: color_data = 12'he61;
			{8'd81, 8'd46}: color_data = 12'he61;
			{8'd81, 8'd47}: color_data = 12'he71;
			{8'd81, 8'd48}: color_data = 12'he71;
			{8'd81, 8'd49}: color_data = 12'he80;
			{8'd81, 8'd50}: color_data = 12'he80;
			{8'd81, 8'd51}: color_data = 12'he80;
			{8'd81, 8'd52}: color_data = 12'he90;
			{8'd81, 8'd53}: color_data = 12'he80;
			{8'd81, 8'd54}: color_data = 12'hff0;
			{8'd81, 8'd125}: color_data = 12'h222;
			{8'd81, 8'd126}: color_data = 12'h111;
			{8'd81, 8'd127}: color_data = 12'h000;
			{8'd81, 8'd128}: color_data = 12'h000;
			{8'd81, 8'd129}: color_data = 12'h000;
			{8'd81, 8'd130}: color_data = 12'h222;
			{8'd81, 8'd131}: color_data = 12'h555;
			{8'd81, 8'd132}: color_data = 12'h777;
			{8'd81, 8'd133}: color_data = 12'h777;
			{8'd81, 8'd134}: color_data = 12'h666;
			{8'd82, 8'd32}: color_data = 12'ha01;
			{8'd82, 8'd33}: color_data = 12'hc01;
			{8'd82, 8'd34}: color_data = 12'hd01;
			{8'd82, 8'd35}: color_data = 12'hd11;
			{8'd82, 8'd36}: color_data = 12'he21;
			{8'd82, 8'd37}: color_data = 12'he21;
			{8'd82, 8'd38}: color_data = 12'he31;
			{8'd82, 8'd39}: color_data = 12'he41;
			{8'd82, 8'd40}: color_data = 12'he41;
			{8'd82, 8'd41}: color_data = 12'he51;
			{8'd82, 8'd42}: color_data = 12'he51;
			{8'd82, 8'd43}: color_data = 12'he51;
			{8'd82, 8'd44}: color_data = 12'he61;
			{8'd82, 8'd45}: color_data = 12'he61;
			{8'd82, 8'd46}: color_data = 12'he61;
			{8'd82, 8'd47}: color_data = 12'he71;
			{8'd82, 8'd48}: color_data = 12'he71;
			{8'd82, 8'd49}: color_data = 12'he80;
			{8'd82, 8'd50}: color_data = 12'he80;
			{8'd82, 8'd51}: color_data = 12'he90;
			{8'd82, 8'd52}: color_data = 12'he90;
			{8'd82, 8'd53}: color_data = 12'he90;
			{8'd82, 8'd54}: color_data = 12'hff0;
			{8'd82, 8'd120}: color_data = 12'h000;
			{8'd82, 8'd121}: color_data = 12'h111;
			{8'd82, 8'd122}: color_data = 12'h111;
			{8'd82, 8'd123}: color_data = 12'h111;
			{8'd82, 8'd124}: color_data = 12'h111;
			{8'd82, 8'd125}: color_data = 12'h111;
			{8'd82, 8'd126}: color_data = 12'h111;
			{8'd82, 8'd127}: color_data = 12'h000;
			{8'd82, 8'd128}: color_data = 12'h222;
			{8'd82, 8'd129}: color_data = 12'h666;
			{8'd82, 8'd130}: color_data = 12'haaa;
			{8'd82, 8'd131}: color_data = 12'hccc;
			{8'd82, 8'd132}: color_data = 12'hbbb;
			{8'd82, 8'd133}: color_data = 12'haaa;
			{8'd82, 8'd134}: color_data = 12'h777;
			{8'd82, 8'd135}: color_data = 12'h444;
			{8'd83, 8'd32}: color_data = 12'hb01;
			{8'd83, 8'd33}: color_data = 12'h901;
			{8'd83, 8'd34}: color_data = 12'h901;
			{8'd83, 8'd35}: color_data = 12'hb11;
			{8'd83, 8'd36}: color_data = 12'hc21;
			{8'd83, 8'd37}: color_data = 12'hd21;
			{8'd83, 8'd38}: color_data = 12'hd31;
			{8'd83, 8'd39}: color_data = 12'hd31;
			{8'd83, 8'd40}: color_data = 12'he41;
			{8'd83, 8'd41}: color_data = 12'he51;
			{8'd83, 8'd42}: color_data = 12'he51;
			{8'd83, 8'd43}: color_data = 12'he51;
			{8'd83, 8'd44}: color_data = 12'he61;
			{8'd83, 8'd45}: color_data = 12'he61;
			{8'd83, 8'd46}: color_data = 12'he61;
			{8'd83, 8'd47}: color_data = 12'he71;
			{8'd83, 8'd48}: color_data = 12'he71;
			{8'd83, 8'd49}: color_data = 12'he80;
			{8'd83, 8'd50}: color_data = 12'he80;
			{8'd83, 8'd51}: color_data = 12'he80;
			{8'd83, 8'd52}: color_data = 12'he90;
			{8'd83, 8'd53}: color_data = 12'hd90;
			{8'd83, 8'd54}: color_data = 12'hff0;
			{8'd83, 8'd114}: color_data = 12'h000;
			{8'd83, 8'd115}: color_data = 12'h222;
			{8'd83, 8'd116}: color_data = 12'h111;
			{8'd83, 8'd117}: color_data = 12'h111;
			{8'd83, 8'd118}: color_data = 12'h111;
			{8'd83, 8'd119}: color_data = 12'h111;
			{8'd83, 8'd120}: color_data = 12'h111;
			{8'd83, 8'd121}: color_data = 12'h111;
			{8'd83, 8'd122}: color_data = 12'h111;
			{8'd83, 8'd123}: color_data = 12'h111;
			{8'd83, 8'd124}: color_data = 12'h111;
			{8'd83, 8'd125}: color_data = 12'h111;
			{8'd83, 8'd126}: color_data = 12'h111;
			{8'd83, 8'd127}: color_data = 12'h111;
			{8'd83, 8'd128}: color_data = 12'h666;
			{8'd83, 8'd129}: color_data = 12'hbbb;
			{8'd83, 8'd130}: color_data = 12'hddd;
			{8'd83, 8'd131}: color_data = 12'heee;
			{8'd83, 8'd132}: color_data = 12'heee;
			{8'd83, 8'd133}: color_data = 12'hddd;
			{8'd83, 8'd134}: color_data = 12'haaa;
			{8'd83, 8'd135}: color_data = 12'h666;
			{8'd83, 8'd136}: color_data = 12'h333;
			{8'd84, 8'd33}: color_data = 12'h700;
			{8'd84, 8'd34}: color_data = 12'h700;
			{8'd84, 8'd35}: color_data = 12'h800;
			{8'd84, 8'd36}: color_data = 12'hb11;
			{8'd84, 8'd37}: color_data = 12'hd21;
			{8'd84, 8'd38}: color_data = 12'hc31;
			{8'd84, 8'd39}: color_data = 12'ha21;
			{8'd84, 8'd40}: color_data = 12'ha31;
			{8'd84, 8'd41}: color_data = 12'hc41;
			{8'd84, 8'd42}: color_data = 12'hd51;
			{8'd84, 8'd43}: color_data = 12'he51;
			{8'd84, 8'd44}: color_data = 12'hd61;
			{8'd84, 8'd45}: color_data = 12'hd61;
			{8'd84, 8'd46}: color_data = 12'he61;
			{8'd84, 8'd47}: color_data = 12'he71;
			{8'd84, 8'd48}: color_data = 12'he71;
			{8'd84, 8'd49}: color_data = 12'he80;
			{8'd84, 8'd50}: color_data = 12'he80;
			{8'd84, 8'd51}: color_data = 12'he80;
			{8'd84, 8'd52}: color_data = 12'he90;
			{8'd84, 8'd53}: color_data = 12'hd80;
			{8'd84, 8'd54}: color_data = 12'hff0;
			{8'd84, 8'd109}: color_data = 12'h000;
			{8'd84, 8'd110}: color_data = 12'h000;
			{8'd84, 8'd111}: color_data = 12'h222;
			{8'd84, 8'd112}: color_data = 12'h222;
			{8'd84, 8'd113}: color_data = 12'h222;
			{8'd84, 8'd114}: color_data = 12'h222;
			{8'd84, 8'd115}: color_data = 12'h222;
			{8'd84, 8'd116}: color_data = 12'h111;
			{8'd84, 8'd117}: color_data = 12'h111;
			{8'd84, 8'd118}: color_data = 12'h111;
			{8'd84, 8'd119}: color_data = 12'h111;
			{8'd84, 8'd120}: color_data = 12'h111;
			{8'd84, 8'd121}: color_data = 12'h111;
			{8'd84, 8'd122}: color_data = 12'h111;
			{8'd84, 8'd123}: color_data = 12'h111;
			{8'd84, 8'd124}: color_data = 12'h111;
			{8'd84, 8'd125}: color_data = 12'h111;
			{8'd84, 8'd126}: color_data = 12'h111;
			{8'd84, 8'd127}: color_data = 12'h333;
			{8'd84, 8'd128}: color_data = 12'h999;
			{8'd84, 8'd129}: color_data = 12'hddd;
			{8'd84, 8'd130}: color_data = 12'hfff;
			{8'd84, 8'd131}: color_data = 12'hfff;
			{8'd84, 8'd132}: color_data = 12'hfff;
			{8'd84, 8'd133}: color_data = 12'heee;
			{8'd84, 8'd134}: color_data = 12'hddd;
			{8'd84, 8'd135}: color_data = 12'h999;
			{8'd84, 8'd136}: color_data = 12'h444;
			{8'd84, 8'd137}: color_data = 12'h222;
			{8'd85, 8'd39}: color_data = 12'h711;
			{8'd85, 8'd40}: color_data = 12'h810;
			{8'd85, 8'd41}: color_data = 12'ha31;
			{8'd85, 8'd42}: color_data = 12'hc41;
			{8'd85, 8'd43}: color_data = 12'he51;
			{8'd85, 8'd44}: color_data = 12'ha41;
			{8'd85, 8'd45}: color_data = 12'h941;
			{8'd85, 8'd46}: color_data = 12'ha50;
			{8'd85, 8'd47}: color_data = 12'hd60;
			{8'd85, 8'd48}: color_data = 12'he70;
			{8'd85, 8'd49}: color_data = 12'hd80;
			{8'd85, 8'd50}: color_data = 12'hd70;
			{8'd85, 8'd51}: color_data = 12'hd80;
			{8'd85, 8'd52}: color_data = 12'he90;
			{8'd85, 8'd53}: color_data = 12'hd80;
			{8'd85, 8'd54}: color_data = 12'h700;
			{8'd85, 8'd104}: color_data = 12'h333;
			{8'd85, 8'd105}: color_data = 12'h222;
			{8'd85, 8'd106}: color_data = 12'h222;
			{8'd85, 8'd107}: color_data = 12'h222;
			{8'd85, 8'd108}: color_data = 12'h222;
			{8'd85, 8'd109}: color_data = 12'h222;
			{8'd85, 8'd110}: color_data = 12'h222;
			{8'd85, 8'd111}: color_data = 12'h222;
			{8'd85, 8'd112}: color_data = 12'h222;
			{8'd85, 8'd113}: color_data = 12'h222;
			{8'd85, 8'd114}: color_data = 12'h222;
			{8'd85, 8'd115}: color_data = 12'h222;
			{8'd85, 8'd116}: color_data = 12'h222;
			{8'd85, 8'd117}: color_data = 12'h111;
			{8'd85, 8'd118}: color_data = 12'h111;
			{8'd85, 8'd119}: color_data = 12'h111;
			{8'd85, 8'd120}: color_data = 12'h111;
			{8'd85, 8'd121}: color_data = 12'h111;
			{8'd85, 8'd122}: color_data = 12'h111;
			{8'd85, 8'd123}: color_data = 12'h111;
			{8'd85, 8'd124}: color_data = 12'h111;
			{8'd85, 8'd125}: color_data = 12'h111;
			{8'd85, 8'd126}: color_data = 12'h111;
			{8'd85, 8'd127}: color_data = 12'h666;
			{8'd85, 8'd128}: color_data = 12'hddd;
			{8'd85, 8'd129}: color_data = 12'hfff;
			{8'd85, 8'd130}: color_data = 12'hfff;
			{8'd85, 8'd131}: color_data = 12'hfff;
			{8'd85, 8'd132}: color_data = 12'hfff;
			{8'd85, 8'd133}: color_data = 12'hfff;
			{8'd85, 8'd134}: color_data = 12'hfff;
			{8'd85, 8'd135}: color_data = 12'hccc;
			{8'd85, 8'd136}: color_data = 12'h777;
			{8'd85, 8'd137}: color_data = 12'h444;
			{8'd86, 8'd45}: color_data = 12'h730;
			{8'd86, 8'd46}: color_data = 12'h830;
			{8'd86, 8'd47}: color_data = 12'hb50;
			{8'd86, 8'd48}: color_data = 12'he70;
			{8'd86, 8'd49}: color_data = 12'hb70;
			{8'd86, 8'd50}: color_data = 12'h950;
			{8'd86, 8'd51}: color_data = 12'h950;
			{8'd86, 8'd52}: color_data = 12'hb70;
			{8'd86, 8'd53}: color_data = 12'hc80;
			{8'd86, 8'd98}: color_data = 12'h000;
			{8'd86, 8'd99}: color_data = 12'h444;
			{8'd86, 8'd100}: color_data = 12'h333;
			{8'd86, 8'd101}: color_data = 12'h333;
			{8'd86, 8'd102}: color_data = 12'h222;
			{8'd86, 8'd103}: color_data = 12'h333;
			{8'd86, 8'd104}: color_data = 12'h222;
			{8'd86, 8'd105}: color_data = 12'h222;
			{8'd86, 8'd106}: color_data = 12'h222;
			{8'd86, 8'd107}: color_data = 12'h222;
			{8'd86, 8'd108}: color_data = 12'h222;
			{8'd86, 8'd109}: color_data = 12'h222;
			{8'd86, 8'd110}: color_data = 12'h222;
			{8'd86, 8'd111}: color_data = 12'h222;
			{8'd86, 8'd112}: color_data = 12'h222;
			{8'd86, 8'd113}: color_data = 12'h222;
			{8'd86, 8'd114}: color_data = 12'h222;
			{8'd86, 8'd115}: color_data = 12'h222;
			{8'd86, 8'd116}: color_data = 12'h222;
			{8'd86, 8'd117}: color_data = 12'h111;
			{8'd86, 8'd118}: color_data = 12'h111;
			{8'd86, 8'd119}: color_data = 12'h111;
			{8'd86, 8'd120}: color_data = 12'h111;
			{8'd86, 8'd121}: color_data = 12'h111;
			{8'd86, 8'd122}: color_data = 12'h111;
			{8'd86, 8'd123}: color_data = 12'h111;
			{8'd86, 8'd124}: color_data = 12'h111;
			{8'd86, 8'd125}: color_data = 12'h111;
			{8'd86, 8'd126}: color_data = 12'h333;
			{8'd86, 8'd127}: color_data = 12'haaa;
			{8'd86, 8'd128}: color_data = 12'heee;
			{8'd86, 8'd129}: color_data = 12'hfff;
			{8'd86, 8'd130}: color_data = 12'hfff;
			{8'd86, 8'd131}: color_data = 12'hfff;
			{8'd86, 8'd132}: color_data = 12'hfff;
			{8'd86, 8'd133}: color_data = 12'hfff;
			{8'd86, 8'd134}: color_data = 12'hfff;
			{8'd86, 8'd135}: color_data = 12'heee;
			{8'd86, 8'd136}: color_data = 12'h999;
			{8'd86, 8'd137}: color_data = 12'h555;
			{8'd87, 8'd50}: color_data = 12'h630;
			{8'd87, 8'd51}: color_data = 12'h740;
			{8'd87, 8'd52}: color_data = 12'h950;
			{8'd87, 8'd53}: color_data = 12'ha70;
			{8'd87, 8'd94}: color_data = 12'h222;
			{8'd87, 8'd95}: color_data = 12'h333;
			{8'd87, 8'd96}: color_data = 12'h333;
			{8'd87, 8'd97}: color_data = 12'h333;
			{8'd87, 8'd98}: color_data = 12'h333;
			{8'd87, 8'd99}: color_data = 12'h333;
			{8'd87, 8'd100}: color_data = 12'h333;
			{8'd87, 8'd101}: color_data = 12'h333;
			{8'd87, 8'd102}: color_data = 12'h333;
			{8'd87, 8'd103}: color_data = 12'h333;
			{8'd87, 8'd104}: color_data = 12'h222;
			{8'd87, 8'd105}: color_data = 12'h222;
			{8'd87, 8'd106}: color_data = 12'h222;
			{8'd87, 8'd107}: color_data = 12'h222;
			{8'd87, 8'd108}: color_data = 12'h222;
			{8'd87, 8'd109}: color_data = 12'h222;
			{8'd87, 8'd110}: color_data = 12'h222;
			{8'd87, 8'd111}: color_data = 12'h222;
			{8'd87, 8'd112}: color_data = 12'h222;
			{8'd87, 8'd113}: color_data = 12'h222;
			{8'd87, 8'd114}: color_data = 12'h222;
			{8'd87, 8'd115}: color_data = 12'h222;
			{8'd87, 8'd116}: color_data = 12'h222;
			{8'd87, 8'd117}: color_data = 12'h222;
			{8'd87, 8'd118}: color_data = 12'h111;
			{8'd87, 8'd119}: color_data = 12'h111;
			{8'd87, 8'd120}: color_data = 12'h111;
			{8'd87, 8'd121}: color_data = 12'h111;
			{8'd87, 8'd122}: color_data = 12'h111;
			{8'd87, 8'd123}: color_data = 12'h111;
			{8'd87, 8'd124}: color_data = 12'h111;
			{8'd87, 8'd125}: color_data = 12'h111;
			{8'd87, 8'd126}: color_data = 12'h555;
			{8'd87, 8'd127}: color_data = 12'hddd;
			{8'd87, 8'd128}: color_data = 12'hfff;
			{8'd87, 8'd129}: color_data = 12'hfff;
			{8'd87, 8'd130}: color_data = 12'hfff;
			{8'd87, 8'd131}: color_data = 12'hfff;
			{8'd87, 8'd132}: color_data = 12'hfff;
			{8'd87, 8'd133}: color_data = 12'hfff;
			{8'd87, 8'd134}: color_data = 12'hfff;
			{8'd87, 8'd135}: color_data = 12'hfff;
			{8'd87, 8'd136}: color_data = 12'hccc;
			{8'd87, 8'd137}: color_data = 12'h777;
			{8'd87, 8'd138}: color_data = 12'h000;
			{8'd88, 8'd88}: color_data = 12'h555;
			{8'd88, 8'd89}: color_data = 12'h444;
			{8'd88, 8'd90}: color_data = 12'h333;
			{8'd88, 8'd91}: color_data = 12'h333;
			{8'd88, 8'd92}: color_data = 12'h333;
			{8'd88, 8'd93}: color_data = 12'h333;
			{8'd88, 8'd94}: color_data = 12'h333;
			{8'd88, 8'd95}: color_data = 12'h333;
			{8'd88, 8'd96}: color_data = 12'h333;
			{8'd88, 8'd97}: color_data = 12'h333;
			{8'd88, 8'd98}: color_data = 12'h333;
			{8'd88, 8'd99}: color_data = 12'h333;
			{8'd88, 8'd100}: color_data = 12'h333;
			{8'd88, 8'd101}: color_data = 12'h333;
			{8'd88, 8'd102}: color_data = 12'h333;
			{8'd88, 8'd103}: color_data = 12'h333;
			{8'd88, 8'd104}: color_data = 12'h222;
			{8'd88, 8'd105}: color_data = 12'h222;
			{8'd88, 8'd106}: color_data = 12'h222;
			{8'd88, 8'd107}: color_data = 12'h222;
			{8'd88, 8'd108}: color_data = 12'h222;
			{8'd88, 8'd109}: color_data = 12'h222;
			{8'd88, 8'd110}: color_data = 12'h222;
			{8'd88, 8'd111}: color_data = 12'h222;
			{8'd88, 8'd112}: color_data = 12'h222;
			{8'd88, 8'd113}: color_data = 12'h222;
			{8'd88, 8'd114}: color_data = 12'h222;
			{8'd88, 8'd115}: color_data = 12'h222;
			{8'd88, 8'd116}: color_data = 12'h222;
			{8'd88, 8'd117}: color_data = 12'h222;
			{8'd88, 8'd118}: color_data = 12'h111;
			{8'd88, 8'd119}: color_data = 12'h111;
			{8'd88, 8'd120}: color_data = 12'h111;
			{8'd88, 8'd121}: color_data = 12'h111;
			{8'd88, 8'd122}: color_data = 12'h111;
			{8'd88, 8'd123}: color_data = 12'h111;
			{8'd88, 8'd124}: color_data = 12'h111;
			{8'd88, 8'd125}: color_data = 12'h222;
			{8'd88, 8'd126}: color_data = 12'h888;
			{8'd88, 8'd127}: color_data = 12'heee;
			{8'd88, 8'd128}: color_data = 12'hfff;
			{8'd88, 8'd129}: color_data = 12'hfff;
			{8'd88, 8'd130}: color_data = 12'hfff;
			{8'd88, 8'd131}: color_data = 12'hfff;
			{8'd88, 8'd132}: color_data = 12'hfff;
			{8'd88, 8'd133}: color_data = 12'hfff;
			{8'd88, 8'd134}: color_data = 12'hfff;
			{8'd88, 8'd135}: color_data = 12'hfff;
			{8'd88, 8'd136}: color_data = 12'heee;
			{8'd88, 8'd137}: color_data = 12'h999;
			{8'd88, 8'd138}: color_data = 12'h555;
			{8'd89, 8'd84}: color_data = 12'h444;
			{8'd89, 8'd85}: color_data = 12'h444;
			{8'd89, 8'd86}: color_data = 12'h444;
			{8'd89, 8'd87}: color_data = 12'h444;
			{8'd89, 8'd88}: color_data = 12'h444;
			{8'd89, 8'd89}: color_data = 12'h444;
			{8'd89, 8'd90}: color_data = 12'h444;
			{8'd89, 8'd91}: color_data = 12'h444;
			{8'd89, 8'd92}: color_data = 12'h333;
			{8'd89, 8'd93}: color_data = 12'h333;
			{8'd89, 8'd94}: color_data = 12'h333;
			{8'd89, 8'd95}: color_data = 12'h333;
			{8'd89, 8'd96}: color_data = 12'h333;
			{8'd89, 8'd97}: color_data = 12'h333;
			{8'd89, 8'd98}: color_data = 12'h333;
			{8'd89, 8'd99}: color_data = 12'h333;
			{8'd89, 8'd100}: color_data = 12'h333;
			{8'd89, 8'd101}: color_data = 12'h333;
			{8'd89, 8'd102}: color_data = 12'h333;
			{8'd89, 8'd103}: color_data = 12'h333;
			{8'd89, 8'd104}: color_data = 12'h222;
			{8'd89, 8'd105}: color_data = 12'h222;
			{8'd89, 8'd106}: color_data = 12'h222;
			{8'd89, 8'd107}: color_data = 12'h222;
			{8'd89, 8'd108}: color_data = 12'h222;
			{8'd89, 8'd109}: color_data = 12'h222;
			{8'd89, 8'd110}: color_data = 12'h222;
			{8'd89, 8'd111}: color_data = 12'h222;
			{8'd89, 8'd112}: color_data = 12'h222;
			{8'd89, 8'd113}: color_data = 12'h222;
			{8'd89, 8'd114}: color_data = 12'h222;
			{8'd89, 8'd115}: color_data = 12'h222;
			{8'd89, 8'd116}: color_data = 12'h222;
			{8'd89, 8'd117}: color_data = 12'h222;
			{8'd89, 8'd118}: color_data = 12'h111;
			{8'd89, 8'd119}: color_data = 12'h111;
			{8'd89, 8'd120}: color_data = 12'h111;
			{8'd89, 8'd121}: color_data = 12'h111;
			{8'd89, 8'd122}: color_data = 12'h111;
			{8'd89, 8'd123}: color_data = 12'h111;
			{8'd89, 8'd124}: color_data = 12'h111;
			{8'd89, 8'd125}: color_data = 12'h333;
			{8'd89, 8'd126}: color_data = 12'hbbb;
			{8'd89, 8'd127}: color_data = 12'hfff;
			{8'd89, 8'd128}: color_data = 12'hfff;
			{8'd89, 8'd129}: color_data = 12'hfff;
			{8'd89, 8'd130}: color_data = 12'hfff;
			{8'd89, 8'd131}: color_data = 12'hfff;
			{8'd89, 8'd132}: color_data = 12'hfff;
			{8'd89, 8'd133}: color_data = 12'hfff;
			{8'd89, 8'd134}: color_data = 12'hfff;
			{8'd89, 8'd135}: color_data = 12'hfff;
			{8'd89, 8'd136}: color_data = 12'hfff;
			{8'd89, 8'd137}: color_data = 12'haaa;
			{8'd89, 8'd138}: color_data = 12'h666;
			{8'd90, 8'd78}: color_data = 12'hfff;
			{8'd90, 8'd79}: color_data = 12'h555;
			{8'd90, 8'd80}: color_data = 12'h444;
			{8'd90, 8'd81}: color_data = 12'h444;
			{8'd90, 8'd82}: color_data = 12'h444;
			{8'd90, 8'd83}: color_data = 12'h444;
			{8'd90, 8'd84}: color_data = 12'h444;
			{8'd90, 8'd85}: color_data = 12'h444;
			{8'd90, 8'd86}: color_data = 12'h444;
			{8'd90, 8'd87}: color_data = 12'h444;
			{8'd90, 8'd88}: color_data = 12'h444;
			{8'd90, 8'd89}: color_data = 12'h444;
			{8'd90, 8'd90}: color_data = 12'h444;
			{8'd90, 8'd91}: color_data = 12'h444;
			{8'd90, 8'd92}: color_data = 12'h444;
			{8'd90, 8'd93}: color_data = 12'h333;
			{8'd90, 8'd94}: color_data = 12'h333;
			{8'd90, 8'd95}: color_data = 12'h333;
			{8'd90, 8'd96}: color_data = 12'h333;
			{8'd90, 8'd97}: color_data = 12'h333;
			{8'd90, 8'd98}: color_data = 12'h333;
			{8'd90, 8'd99}: color_data = 12'h333;
			{8'd90, 8'd100}: color_data = 12'h333;
			{8'd90, 8'd101}: color_data = 12'h333;
			{8'd90, 8'd102}: color_data = 12'h333;
			{8'd90, 8'd103}: color_data = 12'h333;
			{8'd90, 8'd104}: color_data = 12'h333;
			{8'd90, 8'd105}: color_data = 12'h333;
			{8'd90, 8'd106}: color_data = 12'h222;
			{8'd90, 8'd107}: color_data = 12'h222;
			{8'd90, 8'd108}: color_data = 12'h222;
			{8'd90, 8'd109}: color_data = 12'h222;
			{8'd90, 8'd110}: color_data = 12'h222;
			{8'd90, 8'd111}: color_data = 12'h222;
			{8'd90, 8'd112}: color_data = 12'h222;
			{8'd90, 8'd113}: color_data = 12'h222;
			{8'd90, 8'd114}: color_data = 12'h222;
			{8'd90, 8'd115}: color_data = 12'h222;
			{8'd90, 8'd116}: color_data = 12'h222;
			{8'd90, 8'd117}: color_data = 12'h222;
			{8'd90, 8'd118}: color_data = 12'h222;
			{8'd90, 8'd119}: color_data = 12'h111;
			{8'd90, 8'd120}: color_data = 12'h111;
			{8'd90, 8'd121}: color_data = 12'h111;
			{8'd90, 8'd122}: color_data = 12'h111;
			{8'd90, 8'd123}: color_data = 12'h111;
			{8'd90, 8'd124}: color_data = 12'h111;
			{8'd90, 8'd125}: color_data = 12'h555;
			{8'd90, 8'd126}: color_data = 12'hddd;
			{8'd90, 8'd127}: color_data = 12'hfff;
			{8'd90, 8'd128}: color_data = 12'hfff;
			{8'd90, 8'd129}: color_data = 12'hfff;
			{8'd90, 8'd130}: color_data = 12'hfff;
			{8'd90, 8'd131}: color_data = 12'hfff;
			{8'd90, 8'd132}: color_data = 12'hfff;
			{8'd90, 8'd133}: color_data = 12'hfff;
			{8'd90, 8'd134}: color_data = 12'hfff;
			{8'd90, 8'd135}: color_data = 12'hfff;
			{8'd90, 8'd136}: color_data = 12'hfff;
			{8'd90, 8'd137}: color_data = 12'hddd;
			{8'd90, 8'd138}: color_data = 12'h777;
			{8'd90, 8'd139}: color_data = 12'h000;
			{8'd91, 8'd32}: color_data = 12'hf00;
			{8'd91, 8'd33}: color_data = 12'h910;
			{8'd91, 8'd34}: color_data = 12'h920;
			{8'd91, 8'd35}: color_data = 12'h721;
			{8'd91, 8'd73}: color_data = 12'h555;
			{8'd91, 8'd74}: color_data = 12'h444;
			{8'd91, 8'd75}: color_data = 12'h555;
			{8'd91, 8'd76}: color_data = 12'h555;
			{8'd91, 8'd77}: color_data = 12'h555;
			{8'd91, 8'd78}: color_data = 12'h555;
			{8'd91, 8'd79}: color_data = 12'h444;
			{8'd91, 8'd80}: color_data = 12'h444;
			{8'd91, 8'd81}: color_data = 12'h444;
			{8'd91, 8'd82}: color_data = 12'h444;
			{8'd91, 8'd83}: color_data = 12'h444;
			{8'd91, 8'd84}: color_data = 12'h444;
			{8'd91, 8'd85}: color_data = 12'h444;
			{8'd91, 8'd86}: color_data = 12'h444;
			{8'd91, 8'd87}: color_data = 12'h444;
			{8'd91, 8'd88}: color_data = 12'h444;
			{8'd91, 8'd89}: color_data = 12'h444;
			{8'd91, 8'd90}: color_data = 12'h444;
			{8'd91, 8'd91}: color_data = 12'h444;
			{8'd91, 8'd92}: color_data = 12'h333;
			{8'd91, 8'd93}: color_data = 12'h333;
			{8'd91, 8'd94}: color_data = 12'h333;
			{8'd91, 8'd95}: color_data = 12'h333;
			{8'd91, 8'd96}: color_data = 12'h333;
			{8'd91, 8'd97}: color_data = 12'h333;
			{8'd91, 8'd98}: color_data = 12'h333;
			{8'd91, 8'd99}: color_data = 12'h333;
			{8'd91, 8'd100}: color_data = 12'h333;
			{8'd91, 8'd101}: color_data = 12'h333;
			{8'd91, 8'd102}: color_data = 12'h333;
			{8'd91, 8'd103}: color_data = 12'h333;
			{8'd91, 8'd104}: color_data = 12'h333;
			{8'd91, 8'd105}: color_data = 12'h333;
			{8'd91, 8'd106}: color_data = 12'h222;
			{8'd91, 8'd107}: color_data = 12'h222;
			{8'd91, 8'd108}: color_data = 12'h222;
			{8'd91, 8'd109}: color_data = 12'h222;
			{8'd91, 8'd110}: color_data = 12'h222;
			{8'd91, 8'd111}: color_data = 12'h222;
			{8'd91, 8'd112}: color_data = 12'h222;
			{8'd91, 8'd113}: color_data = 12'h222;
			{8'd91, 8'd114}: color_data = 12'h222;
			{8'd91, 8'd115}: color_data = 12'h222;
			{8'd91, 8'd116}: color_data = 12'h222;
			{8'd91, 8'd117}: color_data = 12'h222;
			{8'd91, 8'd118}: color_data = 12'h222;
			{8'd91, 8'd119}: color_data = 12'h222;
			{8'd91, 8'd120}: color_data = 12'h111;
			{8'd91, 8'd121}: color_data = 12'h111;
			{8'd91, 8'd122}: color_data = 12'h111;
			{8'd91, 8'd123}: color_data = 12'h111;
			{8'd91, 8'd124}: color_data = 12'h111;
			{8'd91, 8'd125}: color_data = 12'h888;
			{8'd91, 8'd126}: color_data = 12'heee;
			{8'd91, 8'd127}: color_data = 12'hfff;
			{8'd91, 8'd128}: color_data = 12'hfff;
			{8'd91, 8'd129}: color_data = 12'hfff;
			{8'd91, 8'd130}: color_data = 12'hfff;
			{8'd91, 8'd131}: color_data = 12'hfff;
			{8'd91, 8'd132}: color_data = 12'hfff;
			{8'd91, 8'd133}: color_data = 12'hfff;
			{8'd91, 8'd134}: color_data = 12'hfff;
			{8'd91, 8'd135}: color_data = 12'hfff;
			{8'd91, 8'd136}: color_data = 12'hfff;
			{8'd91, 8'd137}: color_data = 12'heee;
			{8'd91, 8'd138}: color_data = 12'h999;
			{8'd91, 8'd139}: color_data = 12'h444;
			{8'd92, 8'd32}: color_data = 12'ha20;
			{8'd92, 8'd33}: color_data = 12'ha20;
			{8'd92, 8'd34}: color_data = 12'ha21;
			{8'd92, 8'd35}: color_data = 12'ha30;
			{8'd92, 8'd36}: color_data = 12'ha31;
			{8'd92, 8'd37}: color_data = 12'ha30;
			{8'd92, 8'd68}: color_data = 12'h333;
			{8'd92, 8'd69}: color_data = 12'h666;
			{8'd92, 8'd70}: color_data = 12'h555;
			{8'd92, 8'd71}: color_data = 12'h555;
			{8'd92, 8'd72}: color_data = 12'h555;
			{8'd92, 8'd73}: color_data = 12'h555;
			{8'd92, 8'd74}: color_data = 12'h555;
			{8'd92, 8'd75}: color_data = 12'h555;
			{8'd92, 8'd76}: color_data = 12'h555;
			{8'd92, 8'd77}: color_data = 12'h555;
			{8'd92, 8'd78}: color_data = 12'h555;
			{8'd92, 8'd79}: color_data = 12'h555;
			{8'd92, 8'd80}: color_data = 12'h555;
			{8'd92, 8'd81}: color_data = 12'h444;
			{8'd92, 8'd82}: color_data = 12'h444;
			{8'd92, 8'd83}: color_data = 12'h444;
			{8'd92, 8'd84}: color_data = 12'h444;
			{8'd92, 8'd85}: color_data = 12'h444;
			{8'd92, 8'd86}: color_data = 12'h444;
			{8'd92, 8'd87}: color_data = 12'h444;
			{8'd92, 8'd88}: color_data = 12'h444;
			{8'd92, 8'd89}: color_data = 12'h444;
			{8'd92, 8'd90}: color_data = 12'h444;
			{8'd92, 8'd91}: color_data = 12'h444;
			{8'd92, 8'd92}: color_data = 12'h444;
			{8'd92, 8'd93}: color_data = 12'h333;
			{8'd92, 8'd94}: color_data = 12'h333;
			{8'd92, 8'd95}: color_data = 12'h333;
			{8'd92, 8'd96}: color_data = 12'h333;
			{8'd92, 8'd97}: color_data = 12'h333;
			{8'd92, 8'd98}: color_data = 12'h333;
			{8'd92, 8'd99}: color_data = 12'h333;
			{8'd92, 8'd100}: color_data = 12'h333;
			{8'd92, 8'd101}: color_data = 12'h333;
			{8'd92, 8'd102}: color_data = 12'h333;
			{8'd92, 8'd103}: color_data = 12'h333;
			{8'd92, 8'd104}: color_data = 12'h333;
			{8'd92, 8'd105}: color_data = 12'h333;
			{8'd92, 8'd106}: color_data = 12'h333;
			{8'd92, 8'd107}: color_data = 12'h222;
			{8'd92, 8'd108}: color_data = 12'h222;
			{8'd92, 8'd109}: color_data = 12'h222;
			{8'd92, 8'd110}: color_data = 12'h222;
			{8'd92, 8'd111}: color_data = 12'h222;
			{8'd92, 8'd112}: color_data = 12'h222;
			{8'd92, 8'd113}: color_data = 12'h222;
			{8'd92, 8'd114}: color_data = 12'h222;
			{8'd92, 8'd115}: color_data = 12'h222;
			{8'd92, 8'd116}: color_data = 12'h222;
			{8'd92, 8'd117}: color_data = 12'h222;
			{8'd92, 8'd118}: color_data = 12'h222;
			{8'd92, 8'd119}: color_data = 12'h222;
			{8'd92, 8'd120}: color_data = 12'h111;
			{8'd92, 8'd121}: color_data = 12'h111;
			{8'd92, 8'd122}: color_data = 12'h111;
			{8'd92, 8'd123}: color_data = 12'h111;
			{8'd92, 8'd124}: color_data = 12'h222;
			{8'd92, 8'd125}: color_data = 12'haaa;
			{8'd92, 8'd126}: color_data = 12'hfff;
			{8'd92, 8'd127}: color_data = 12'hfff;
			{8'd92, 8'd128}: color_data = 12'hfff;
			{8'd92, 8'd129}: color_data = 12'hfff;
			{8'd92, 8'd130}: color_data = 12'hfff;
			{8'd92, 8'd131}: color_data = 12'hfff;
			{8'd92, 8'd132}: color_data = 12'hfff;
			{8'd92, 8'd133}: color_data = 12'hfff;
			{8'd92, 8'd134}: color_data = 12'hfff;
			{8'd92, 8'd135}: color_data = 12'hfff;
			{8'd92, 8'd136}: color_data = 12'hfff;
			{8'd92, 8'd137}: color_data = 12'hfff;
			{8'd92, 8'd138}: color_data = 12'haaa;
			{8'd92, 8'd139}: color_data = 12'h777;
			{8'd93, 8'd32}: color_data = 12'ha20;
			{8'd93, 8'd33}: color_data = 12'hc21;
			{8'd93, 8'd34}: color_data = 12'hd31;
			{8'd93, 8'd35}: color_data = 12'hd41;
			{8'd93, 8'd36}: color_data = 12'hd41;
			{8'd93, 8'd37}: color_data = 12'hb41;
			{8'd93, 8'd38}: color_data = 12'ha30;
			{8'd93, 8'd39}: color_data = 12'ha40;
			{8'd93, 8'd40}: color_data = 12'ha40;
			{8'd93, 8'd41}: color_data = 12'ha50;
			{8'd93, 8'd42}: color_data = 12'ha50;
			{8'd93, 8'd43}: color_data = 12'ha50;
			{8'd93, 8'd44}: color_data = 12'ha50;
			{8'd93, 8'd45}: color_data = 12'ha60;
			{8'd93, 8'd46}: color_data = 12'ha60;
			{8'd93, 8'd47}: color_data = 12'ha60;
			{8'd93, 8'd48}: color_data = 12'ha60;
			{8'd93, 8'd49}: color_data = 12'ha60;
			{8'd93, 8'd50}: color_data = 12'ha70;
			{8'd93, 8'd51}: color_data = 12'h970;
			{8'd93, 8'd52}: color_data = 12'h960;
			{8'd93, 8'd63}: color_data = 12'h666;
			{8'd93, 8'd64}: color_data = 12'h555;
			{8'd93, 8'd65}: color_data = 12'h666;
			{8'd93, 8'd66}: color_data = 12'h555;
			{8'd93, 8'd67}: color_data = 12'h555;
			{8'd93, 8'd68}: color_data = 12'h555;
			{8'd93, 8'd69}: color_data = 12'h555;
			{8'd93, 8'd70}: color_data = 12'h555;
			{8'd93, 8'd71}: color_data = 12'h555;
			{8'd93, 8'd72}: color_data = 12'h555;
			{8'd93, 8'd73}: color_data = 12'h555;
			{8'd93, 8'd74}: color_data = 12'h555;
			{8'd93, 8'd75}: color_data = 12'h555;
			{8'd93, 8'd76}: color_data = 12'h555;
			{8'd93, 8'd77}: color_data = 12'h555;
			{8'd93, 8'd78}: color_data = 12'h555;
			{8'd93, 8'd79}: color_data = 12'h555;
			{8'd93, 8'd80}: color_data = 12'h444;
			{8'd93, 8'd81}: color_data = 12'h444;
			{8'd93, 8'd82}: color_data = 12'h444;
			{8'd93, 8'd83}: color_data = 12'h444;
			{8'd93, 8'd84}: color_data = 12'h444;
			{8'd93, 8'd85}: color_data = 12'h444;
			{8'd93, 8'd86}: color_data = 12'h444;
			{8'd93, 8'd87}: color_data = 12'h444;
			{8'd93, 8'd88}: color_data = 12'h444;
			{8'd93, 8'd89}: color_data = 12'h444;
			{8'd93, 8'd90}: color_data = 12'h444;
			{8'd93, 8'd91}: color_data = 12'h444;
			{8'd93, 8'd92}: color_data = 12'h444;
			{8'd93, 8'd93}: color_data = 12'h444;
			{8'd93, 8'd94}: color_data = 12'h333;
			{8'd93, 8'd95}: color_data = 12'h333;
			{8'd93, 8'd96}: color_data = 12'h333;
			{8'd93, 8'd97}: color_data = 12'h333;
			{8'd93, 8'd98}: color_data = 12'h333;
			{8'd93, 8'd99}: color_data = 12'h333;
			{8'd93, 8'd100}: color_data = 12'h333;
			{8'd93, 8'd101}: color_data = 12'h333;
			{8'd93, 8'd102}: color_data = 12'h333;
			{8'd93, 8'd103}: color_data = 12'h333;
			{8'd93, 8'd104}: color_data = 12'h333;
			{8'd93, 8'd105}: color_data = 12'h333;
			{8'd93, 8'd106}: color_data = 12'h333;
			{8'd93, 8'd107}: color_data = 12'h222;
			{8'd93, 8'd108}: color_data = 12'h222;
			{8'd93, 8'd109}: color_data = 12'h222;
			{8'd93, 8'd110}: color_data = 12'h222;
			{8'd93, 8'd111}: color_data = 12'h222;
			{8'd93, 8'd112}: color_data = 12'h222;
			{8'd93, 8'd113}: color_data = 12'h222;
			{8'd93, 8'd114}: color_data = 12'h222;
			{8'd93, 8'd115}: color_data = 12'h222;
			{8'd93, 8'd116}: color_data = 12'h222;
			{8'd93, 8'd117}: color_data = 12'h222;
			{8'd93, 8'd118}: color_data = 12'h222;
			{8'd93, 8'd119}: color_data = 12'h222;
			{8'd93, 8'd120}: color_data = 12'h111;
			{8'd93, 8'd121}: color_data = 12'h111;
			{8'd93, 8'd122}: color_data = 12'h111;
			{8'd93, 8'd123}: color_data = 12'h111;
			{8'd93, 8'd124}: color_data = 12'h333;
			{8'd93, 8'd125}: color_data = 12'hccc;
			{8'd93, 8'd126}: color_data = 12'hfff;
			{8'd93, 8'd127}: color_data = 12'hfff;
			{8'd93, 8'd128}: color_data = 12'hfff;
			{8'd93, 8'd129}: color_data = 12'hfff;
			{8'd93, 8'd130}: color_data = 12'hfff;
			{8'd93, 8'd131}: color_data = 12'hfff;
			{8'd93, 8'd132}: color_data = 12'hfff;
			{8'd93, 8'd133}: color_data = 12'hfff;
			{8'd93, 8'd134}: color_data = 12'hfff;
			{8'd93, 8'd135}: color_data = 12'hfff;
			{8'd93, 8'd136}: color_data = 12'hfff;
			{8'd93, 8'd137}: color_data = 12'hfff;
			{8'd93, 8'd138}: color_data = 12'hbbb;
			{8'd93, 8'd139}: color_data = 12'h777;
			{8'd94, 8'd32}: color_data = 12'ha21;
			{8'd94, 8'd33}: color_data = 12'hc21;
			{8'd94, 8'd34}: color_data = 12'hd31;
			{8'd94, 8'd35}: color_data = 12'he41;
			{8'd94, 8'd36}: color_data = 12'he41;
			{8'd94, 8'd37}: color_data = 12'hd51;
			{8'd94, 8'd38}: color_data = 12'hc41;
			{8'd94, 8'd39}: color_data = 12'hb51;
			{8'd94, 8'd40}: color_data = 12'hb51;
			{8'd94, 8'd41}: color_data = 12'hb51;
			{8'd94, 8'd42}: color_data = 12'hb61;
			{8'd94, 8'd43}: color_data = 12'hb61;
			{8'd94, 8'd44}: color_data = 12'hb60;
			{8'd94, 8'd45}: color_data = 12'hb60;
			{8'd94, 8'd46}: color_data = 12'hb70;
			{8'd94, 8'd47}: color_data = 12'hb70;
			{8'd94, 8'd48}: color_data = 12'hb70;
			{8'd94, 8'd49}: color_data = 12'hb70;
			{8'd94, 8'd50}: color_data = 12'hb80;
			{8'd94, 8'd51}: color_data = 12'hb80;
			{8'd94, 8'd52}: color_data = 12'ha70;
			{8'd94, 8'd57}: color_data = 12'h555;
			{8'd94, 8'd58}: color_data = 12'h666;
			{8'd94, 8'd59}: color_data = 12'h666;
			{8'd94, 8'd60}: color_data = 12'h666;
			{8'd94, 8'd61}: color_data = 12'h666;
			{8'd94, 8'd62}: color_data = 12'h666;
			{8'd94, 8'd63}: color_data = 12'h666;
			{8'd94, 8'd64}: color_data = 12'h666;
			{8'd94, 8'd65}: color_data = 12'h666;
			{8'd94, 8'd66}: color_data = 12'h666;
			{8'd94, 8'd67}: color_data = 12'h666;
			{8'd94, 8'd68}: color_data = 12'h666;
			{8'd94, 8'd69}: color_data = 12'h555;
			{8'd94, 8'd70}: color_data = 12'h555;
			{8'd94, 8'd71}: color_data = 12'h555;
			{8'd94, 8'd72}: color_data = 12'h555;
			{8'd94, 8'd73}: color_data = 12'h555;
			{8'd94, 8'd74}: color_data = 12'h555;
			{8'd94, 8'd75}: color_data = 12'h555;
			{8'd94, 8'd76}: color_data = 12'h555;
			{8'd94, 8'd77}: color_data = 12'h555;
			{8'd94, 8'd78}: color_data = 12'h555;
			{8'd94, 8'd79}: color_data = 12'h555;
			{8'd94, 8'd80}: color_data = 12'h444;
			{8'd94, 8'd81}: color_data = 12'h444;
			{8'd94, 8'd82}: color_data = 12'h444;
			{8'd94, 8'd83}: color_data = 12'h444;
			{8'd94, 8'd84}: color_data = 12'h444;
			{8'd94, 8'd85}: color_data = 12'h444;
			{8'd94, 8'd86}: color_data = 12'h444;
			{8'd94, 8'd87}: color_data = 12'h444;
			{8'd94, 8'd88}: color_data = 12'h444;
			{8'd94, 8'd89}: color_data = 12'h444;
			{8'd94, 8'd90}: color_data = 12'h444;
			{8'd94, 8'd91}: color_data = 12'h444;
			{8'd94, 8'd92}: color_data = 12'h444;
			{8'd94, 8'd93}: color_data = 12'h444;
			{8'd94, 8'd94}: color_data = 12'h333;
			{8'd94, 8'd95}: color_data = 12'h333;
			{8'd94, 8'd96}: color_data = 12'h333;
			{8'd94, 8'd97}: color_data = 12'h333;
			{8'd94, 8'd98}: color_data = 12'h333;
			{8'd94, 8'd99}: color_data = 12'h333;
			{8'd94, 8'd100}: color_data = 12'h333;
			{8'd94, 8'd101}: color_data = 12'h333;
			{8'd94, 8'd102}: color_data = 12'h333;
			{8'd94, 8'd103}: color_data = 12'h333;
			{8'd94, 8'd104}: color_data = 12'h333;
			{8'd94, 8'd105}: color_data = 12'h333;
			{8'd94, 8'd106}: color_data = 12'h333;
			{8'd94, 8'd107}: color_data = 12'h222;
			{8'd94, 8'd108}: color_data = 12'h222;
			{8'd94, 8'd109}: color_data = 12'h222;
			{8'd94, 8'd110}: color_data = 12'h222;
			{8'd94, 8'd111}: color_data = 12'h222;
			{8'd94, 8'd112}: color_data = 12'h222;
			{8'd94, 8'd113}: color_data = 12'h222;
			{8'd94, 8'd114}: color_data = 12'h222;
			{8'd94, 8'd115}: color_data = 12'h222;
			{8'd94, 8'd116}: color_data = 12'h222;
			{8'd94, 8'd117}: color_data = 12'h222;
			{8'd94, 8'd118}: color_data = 12'h222;
			{8'd94, 8'd119}: color_data = 12'h222;
			{8'd94, 8'd120}: color_data = 12'h111;
			{8'd94, 8'd121}: color_data = 12'h111;
			{8'd94, 8'd122}: color_data = 12'h111;
			{8'd94, 8'd123}: color_data = 12'h111;
			{8'd94, 8'd124}: color_data = 12'h555;
			{8'd94, 8'd125}: color_data = 12'heee;
			{8'd94, 8'd126}: color_data = 12'hfff;
			{8'd94, 8'd127}: color_data = 12'hfff;
			{8'd94, 8'd128}: color_data = 12'hfff;
			{8'd94, 8'd129}: color_data = 12'hfff;
			{8'd94, 8'd130}: color_data = 12'hfff;
			{8'd94, 8'd131}: color_data = 12'hfff;
			{8'd94, 8'd132}: color_data = 12'hfff;
			{8'd94, 8'd133}: color_data = 12'hfff;
			{8'd94, 8'd134}: color_data = 12'hfff;
			{8'd94, 8'd135}: color_data = 12'hfff;
			{8'd94, 8'd136}: color_data = 12'hfff;
			{8'd94, 8'd137}: color_data = 12'hfff;
			{8'd94, 8'd138}: color_data = 12'hddd;
			{8'd94, 8'd139}: color_data = 12'h777;
			{8'd94, 8'd140}: color_data = 12'h000;
			{8'd95, 8'd32}: color_data = 12'h920;
			{8'd95, 8'd33}: color_data = 12'hc21;
			{8'd95, 8'd34}: color_data = 12'he31;
			{8'd95, 8'd35}: color_data = 12'he41;
			{8'd95, 8'd36}: color_data = 12'he41;
			{8'd95, 8'd37}: color_data = 12'he51;
			{8'd95, 8'd38}: color_data = 12'he51;
			{8'd95, 8'd39}: color_data = 12'he61;
			{8'd95, 8'd40}: color_data = 12'he61;
			{8'd95, 8'd41}: color_data = 12'he61;
			{8'd95, 8'd42}: color_data = 12'he71;
			{8'd95, 8'd43}: color_data = 12'he71;
			{8'd95, 8'd44}: color_data = 12'he71;
			{8'd95, 8'd45}: color_data = 12'he80;
			{8'd95, 8'd46}: color_data = 12'he80;
			{8'd95, 8'd47}: color_data = 12'he80;
			{8'd95, 8'd48}: color_data = 12'he90;
			{8'd95, 8'd49}: color_data = 12'he90;
			{8'd95, 8'd50}: color_data = 12'he90;
			{8'd95, 8'd51}: color_data = 12'he90;
			{8'd95, 8'd52}: color_data = 12'hc80;
			{8'd95, 8'd54}: color_data = 12'h777;
			{8'd95, 8'd55}: color_data = 12'h666;
			{8'd95, 8'd56}: color_data = 12'h666;
			{8'd95, 8'd57}: color_data = 12'h666;
			{8'd95, 8'd58}: color_data = 12'h666;
			{8'd95, 8'd59}: color_data = 12'h666;
			{8'd95, 8'd60}: color_data = 12'h666;
			{8'd95, 8'd61}: color_data = 12'h666;
			{8'd95, 8'd62}: color_data = 12'h666;
			{8'd95, 8'd63}: color_data = 12'h666;
			{8'd95, 8'd64}: color_data = 12'h666;
			{8'd95, 8'd65}: color_data = 12'h666;
			{8'd95, 8'd66}: color_data = 12'h666;
			{8'd95, 8'd67}: color_data = 12'h666;
			{8'd95, 8'd68}: color_data = 12'h555;
			{8'd95, 8'd69}: color_data = 12'h555;
			{8'd95, 8'd70}: color_data = 12'h555;
			{8'd95, 8'd71}: color_data = 12'h555;
			{8'd95, 8'd72}: color_data = 12'h555;
			{8'd95, 8'd73}: color_data = 12'h555;
			{8'd95, 8'd74}: color_data = 12'h555;
			{8'd95, 8'd75}: color_data = 12'h555;
			{8'd95, 8'd76}: color_data = 12'h555;
			{8'd95, 8'd77}: color_data = 12'h555;
			{8'd95, 8'd78}: color_data = 12'h555;
			{8'd95, 8'd79}: color_data = 12'h555;
			{8'd95, 8'd80}: color_data = 12'h444;
			{8'd95, 8'd81}: color_data = 12'h444;
			{8'd95, 8'd82}: color_data = 12'h444;
			{8'd95, 8'd83}: color_data = 12'h444;
			{8'd95, 8'd84}: color_data = 12'h444;
			{8'd95, 8'd85}: color_data = 12'h444;
			{8'd95, 8'd86}: color_data = 12'h444;
			{8'd95, 8'd87}: color_data = 12'h444;
			{8'd95, 8'd88}: color_data = 12'h444;
			{8'd95, 8'd89}: color_data = 12'h444;
			{8'd95, 8'd90}: color_data = 12'h444;
			{8'd95, 8'd91}: color_data = 12'h444;
			{8'd95, 8'd92}: color_data = 12'h444;
			{8'd95, 8'd93}: color_data = 12'h444;
			{8'd95, 8'd94}: color_data = 12'h333;
			{8'd95, 8'd95}: color_data = 12'h333;
			{8'd95, 8'd96}: color_data = 12'h333;
			{8'd95, 8'd97}: color_data = 12'h333;
			{8'd95, 8'd98}: color_data = 12'h333;
			{8'd95, 8'd99}: color_data = 12'h333;
			{8'd95, 8'd100}: color_data = 12'h333;
			{8'd95, 8'd101}: color_data = 12'h333;
			{8'd95, 8'd102}: color_data = 12'h333;
			{8'd95, 8'd103}: color_data = 12'h333;
			{8'd95, 8'd104}: color_data = 12'h333;
			{8'd95, 8'd105}: color_data = 12'h333;
			{8'd95, 8'd106}: color_data = 12'h333;
			{8'd95, 8'd107}: color_data = 12'h222;
			{8'd95, 8'd108}: color_data = 12'h222;
			{8'd95, 8'd109}: color_data = 12'h222;
			{8'd95, 8'd110}: color_data = 12'h222;
			{8'd95, 8'd111}: color_data = 12'h222;
			{8'd95, 8'd112}: color_data = 12'h222;
			{8'd95, 8'd113}: color_data = 12'h222;
			{8'd95, 8'd114}: color_data = 12'h222;
			{8'd95, 8'd115}: color_data = 12'h222;
			{8'd95, 8'd116}: color_data = 12'h222;
			{8'd95, 8'd117}: color_data = 12'h222;
			{8'd95, 8'd118}: color_data = 12'h222;
			{8'd95, 8'd119}: color_data = 12'h222;
			{8'd95, 8'd120}: color_data = 12'h222;
			{8'd95, 8'd121}: color_data = 12'h111;
			{8'd95, 8'd122}: color_data = 12'h111;
			{8'd95, 8'd123}: color_data = 12'h111;
			{8'd95, 8'd124}: color_data = 12'h777;
			{8'd95, 8'd125}: color_data = 12'hfff;
			{8'd95, 8'd126}: color_data = 12'hfff;
			{8'd95, 8'd127}: color_data = 12'hfff;
			{8'd95, 8'd128}: color_data = 12'hfff;
			{8'd95, 8'd129}: color_data = 12'hfff;
			{8'd95, 8'd130}: color_data = 12'hfff;
			{8'd95, 8'd131}: color_data = 12'hfff;
			{8'd95, 8'd132}: color_data = 12'hfff;
			{8'd95, 8'd133}: color_data = 12'hfff;
			{8'd95, 8'd134}: color_data = 12'hfff;
			{8'd95, 8'd135}: color_data = 12'hfff;
			{8'd95, 8'd136}: color_data = 12'hfff;
			{8'd95, 8'd137}: color_data = 12'hfff;
			{8'd95, 8'd138}: color_data = 12'heee;
			{8'd95, 8'd139}: color_data = 12'h999;
			{8'd95, 8'd140}: color_data = 12'h222;
			{8'd96, 8'd32}: color_data = 12'hd21;
			{8'd96, 8'd33}: color_data = 12'hd31;
			{8'd96, 8'd34}: color_data = 12'he31;
			{8'd96, 8'd35}: color_data = 12'he41;
			{8'd96, 8'd36}: color_data = 12'he41;
			{8'd96, 8'd37}: color_data = 12'he51;
			{8'd96, 8'd38}: color_data = 12'he51;
			{8'd96, 8'd39}: color_data = 12'he51;
			{8'd96, 8'd40}: color_data = 12'he61;
			{8'd96, 8'd41}: color_data = 12'he61;
			{8'd96, 8'd42}: color_data = 12'he71;
			{8'd96, 8'd43}: color_data = 12'he71;
			{8'd96, 8'd44}: color_data = 12'he71;
			{8'd96, 8'd45}: color_data = 12'he80;
			{8'd96, 8'd46}: color_data = 12'he80;
			{8'd96, 8'd47}: color_data = 12'he80;
			{8'd96, 8'd48}: color_data = 12'he90;
			{8'd96, 8'd49}: color_data = 12'he90;
			{8'd96, 8'd50}: color_data = 12'he90;
			{8'd96, 8'd51}: color_data = 12'hea0;
			{8'd96, 8'd52}: color_data = 12'hea0;
			{8'd96, 8'd53}: color_data = 12'h35a;
			{8'd96, 8'd54}: color_data = 12'h666;
			{8'd96, 8'd55}: color_data = 12'h666;
			{8'd96, 8'd56}: color_data = 12'h666;
			{8'd96, 8'd57}: color_data = 12'h666;
			{8'd96, 8'd58}: color_data = 12'h666;
			{8'd96, 8'd59}: color_data = 12'h666;
			{8'd96, 8'd60}: color_data = 12'h666;
			{8'd96, 8'd61}: color_data = 12'h666;
			{8'd96, 8'd62}: color_data = 12'h666;
			{8'd96, 8'd63}: color_data = 12'h666;
			{8'd96, 8'd64}: color_data = 12'h666;
			{8'd96, 8'd65}: color_data = 12'h666;
			{8'd96, 8'd66}: color_data = 12'h666;
			{8'd96, 8'd67}: color_data = 12'h666;
			{8'd96, 8'd68}: color_data = 12'h555;
			{8'd96, 8'd69}: color_data = 12'h555;
			{8'd96, 8'd70}: color_data = 12'h555;
			{8'd96, 8'd71}: color_data = 12'h555;
			{8'd96, 8'd72}: color_data = 12'h555;
			{8'd96, 8'd73}: color_data = 12'h555;
			{8'd96, 8'd74}: color_data = 12'h555;
			{8'd96, 8'd75}: color_data = 12'h555;
			{8'd96, 8'd76}: color_data = 12'h555;
			{8'd96, 8'd77}: color_data = 12'h555;
			{8'd96, 8'd78}: color_data = 12'h555;
			{8'd96, 8'd79}: color_data = 12'h555;
			{8'd96, 8'd80}: color_data = 12'h555;
			{8'd96, 8'd81}: color_data = 12'h444;
			{8'd96, 8'd82}: color_data = 12'h444;
			{8'd96, 8'd83}: color_data = 12'h444;
			{8'd96, 8'd84}: color_data = 12'h444;
			{8'd96, 8'd85}: color_data = 12'h444;
			{8'd96, 8'd86}: color_data = 12'h444;
			{8'd96, 8'd87}: color_data = 12'h444;
			{8'd96, 8'd88}: color_data = 12'h444;
			{8'd96, 8'd89}: color_data = 12'h444;
			{8'd96, 8'd90}: color_data = 12'h444;
			{8'd96, 8'd91}: color_data = 12'h444;
			{8'd96, 8'd92}: color_data = 12'h444;
			{8'd96, 8'd93}: color_data = 12'h444;
			{8'd96, 8'd94}: color_data = 12'h333;
			{8'd96, 8'd95}: color_data = 12'h333;
			{8'd96, 8'd96}: color_data = 12'h333;
			{8'd96, 8'd97}: color_data = 12'h333;
			{8'd96, 8'd98}: color_data = 12'h333;
			{8'd96, 8'd99}: color_data = 12'h333;
			{8'd96, 8'd100}: color_data = 12'h333;
			{8'd96, 8'd101}: color_data = 12'h333;
			{8'd96, 8'd102}: color_data = 12'h333;
			{8'd96, 8'd103}: color_data = 12'h333;
			{8'd96, 8'd104}: color_data = 12'h333;
			{8'd96, 8'd105}: color_data = 12'h333;
			{8'd96, 8'd106}: color_data = 12'h333;
			{8'd96, 8'd107}: color_data = 12'h222;
			{8'd96, 8'd108}: color_data = 12'h222;
			{8'd96, 8'd109}: color_data = 12'h222;
			{8'd96, 8'd110}: color_data = 12'h222;
			{8'd96, 8'd111}: color_data = 12'h222;
			{8'd96, 8'd112}: color_data = 12'h222;
			{8'd96, 8'd113}: color_data = 12'h222;
			{8'd96, 8'd114}: color_data = 12'h222;
			{8'd96, 8'd115}: color_data = 12'h222;
			{8'd96, 8'd116}: color_data = 12'h222;
			{8'd96, 8'd117}: color_data = 12'h222;
			{8'd96, 8'd118}: color_data = 12'h222;
			{8'd96, 8'd119}: color_data = 12'h222;
			{8'd96, 8'd120}: color_data = 12'h222;
			{8'd96, 8'd121}: color_data = 12'h111;
			{8'd96, 8'd122}: color_data = 12'h111;
			{8'd96, 8'd123}: color_data = 12'h111;
			{8'd96, 8'd124}: color_data = 12'h999;
			{8'd96, 8'd125}: color_data = 12'hfff;
			{8'd96, 8'd126}: color_data = 12'hfff;
			{8'd96, 8'd127}: color_data = 12'hfff;
			{8'd96, 8'd128}: color_data = 12'hfff;
			{8'd96, 8'd129}: color_data = 12'hfff;
			{8'd96, 8'd130}: color_data = 12'hfff;
			{8'd96, 8'd131}: color_data = 12'hfff;
			{8'd96, 8'd132}: color_data = 12'hfff;
			{8'd96, 8'd133}: color_data = 12'hfff;
			{8'd96, 8'd134}: color_data = 12'hfff;
			{8'd96, 8'd135}: color_data = 12'hfff;
			{8'd96, 8'd136}: color_data = 12'hfff;
			{8'd96, 8'd137}: color_data = 12'hfff;
			{8'd96, 8'd138}: color_data = 12'heee;
			{8'd96, 8'd139}: color_data = 12'h999;
			{8'd96, 8'd140}: color_data = 12'h555;
			{8'd97, 8'd32}: color_data = 12'hc21;
			{8'd97, 8'd33}: color_data = 12'hd31;
			{8'd97, 8'd34}: color_data = 12'he31;
			{8'd97, 8'd35}: color_data = 12'he41;
			{8'd97, 8'd36}: color_data = 12'he41;
			{8'd97, 8'd37}: color_data = 12'he51;
			{8'd97, 8'd38}: color_data = 12'he51;
			{8'd97, 8'd39}: color_data = 12'he51;
			{8'd97, 8'd40}: color_data = 12'he61;
			{8'd97, 8'd41}: color_data = 12'he61;
			{8'd97, 8'd42}: color_data = 12'he71;
			{8'd97, 8'd43}: color_data = 12'he71;
			{8'd97, 8'd44}: color_data = 12'he71;
			{8'd97, 8'd45}: color_data = 12'he80;
			{8'd97, 8'd46}: color_data = 12'he80;
			{8'd97, 8'd47}: color_data = 12'he80;
			{8'd97, 8'd48}: color_data = 12'he90;
			{8'd97, 8'd49}: color_data = 12'he90;
			{8'd97, 8'd50}: color_data = 12'he90;
			{8'd97, 8'd51}: color_data = 12'hea0;
			{8'd97, 8'd52}: color_data = 12'hea0;
			{8'd97, 8'd53}: color_data = 12'h458;
			{8'd97, 8'd54}: color_data = 12'h777;
			{8'd97, 8'd55}: color_data = 12'h777;
			{8'd97, 8'd56}: color_data = 12'h666;
			{8'd97, 8'd57}: color_data = 12'h666;
			{8'd97, 8'd58}: color_data = 12'h666;
			{8'd97, 8'd59}: color_data = 12'h666;
			{8'd97, 8'd60}: color_data = 12'h666;
			{8'd97, 8'd61}: color_data = 12'h666;
			{8'd97, 8'd62}: color_data = 12'h666;
			{8'd97, 8'd63}: color_data = 12'h666;
			{8'd97, 8'd64}: color_data = 12'h666;
			{8'd97, 8'd65}: color_data = 12'h666;
			{8'd97, 8'd66}: color_data = 12'h666;
			{8'd97, 8'd67}: color_data = 12'h666;
			{8'd97, 8'd68}: color_data = 12'h555;
			{8'd97, 8'd69}: color_data = 12'h555;
			{8'd97, 8'd70}: color_data = 12'h555;
			{8'd97, 8'd71}: color_data = 12'h555;
			{8'd97, 8'd72}: color_data = 12'h555;
			{8'd97, 8'd73}: color_data = 12'h555;
			{8'd97, 8'd74}: color_data = 12'h555;
			{8'd97, 8'd75}: color_data = 12'h555;
			{8'd97, 8'd76}: color_data = 12'h555;
			{8'd97, 8'd77}: color_data = 12'h555;
			{8'd97, 8'd78}: color_data = 12'h555;
			{8'd97, 8'd79}: color_data = 12'h555;
			{8'd97, 8'd80}: color_data = 12'h555;
			{8'd97, 8'd81}: color_data = 12'h444;
			{8'd97, 8'd82}: color_data = 12'h444;
			{8'd97, 8'd83}: color_data = 12'h444;
			{8'd97, 8'd84}: color_data = 12'h444;
			{8'd97, 8'd85}: color_data = 12'h444;
			{8'd97, 8'd86}: color_data = 12'h444;
			{8'd97, 8'd87}: color_data = 12'h444;
			{8'd97, 8'd88}: color_data = 12'h444;
			{8'd97, 8'd89}: color_data = 12'h444;
			{8'd97, 8'd90}: color_data = 12'h444;
			{8'd97, 8'd91}: color_data = 12'h444;
			{8'd97, 8'd92}: color_data = 12'h444;
			{8'd97, 8'd93}: color_data = 12'h444;
			{8'd97, 8'd94}: color_data = 12'h333;
			{8'd97, 8'd95}: color_data = 12'h333;
			{8'd97, 8'd96}: color_data = 12'h333;
			{8'd97, 8'd97}: color_data = 12'h333;
			{8'd97, 8'd98}: color_data = 12'h333;
			{8'd97, 8'd99}: color_data = 12'h333;
			{8'd97, 8'd100}: color_data = 12'h333;
			{8'd97, 8'd101}: color_data = 12'h333;
			{8'd97, 8'd102}: color_data = 12'h333;
			{8'd97, 8'd103}: color_data = 12'h333;
			{8'd97, 8'd104}: color_data = 12'h333;
			{8'd97, 8'd105}: color_data = 12'h333;
			{8'd97, 8'd106}: color_data = 12'h333;
			{8'd97, 8'd107}: color_data = 12'h222;
			{8'd97, 8'd108}: color_data = 12'h222;
			{8'd97, 8'd109}: color_data = 12'h222;
			{8'd97, 8'd110}: color_data = 12'h222;
			{8'd97, 8'd111}: color_data = 12'h222;
			{8'd97, 8'd112}: color_data = 12'h222;
			{8'd97, 8'd113}: color_data = 12'h222;
			{8'd97, 8'd114}: color_data = 12'h222;
			{8'd97, 8'd115}: color_data = 12'h222;
			{8'd97, 8'd116}: color_data = 12'h222;
			{8'd97, 8'd117}: color_data = 12'h222;
			{8'd97, 8'd118}: color_data = 12'h222;
			{8'd97, 8'd119}: color_data = 12'h222;
			{8'd97, 8'd120}: color_data = 12'h222;
			{8'd97, 8'd121}: color_data = 12'h111;
			{8'd97, 8'd122}: color_data = 12'h111;
			{8'd97, 8'd123}: color_data = 12'h222;
			{8'd97, 8'd124}: color_data = 12'hbbb;
			{8'd97, 8'd125}: color_data = 12'hfff;
			{8'd97, 8'd126}: color_data = 12'hfff;
			{8'd97, 8'd127}: color_data = 12'hfff;
			{8'd97, 8'd128}: color_data = 12'hfff;
			{8'd97, 8'd129}: color_data = 12'hfff;
			{8'd97, 8'd130}: color_data = 12'hfff;
			{8'd97, 8'd131}: color_data = 12'hfff;
			{8'd97, 8'd132}: color_data = 12'hfff;
			{8'd97, 8'd133}: color_data = 12'hfff;
			{8'd97, 8'd134}: color_data = 12'hfff;
			{8'd97, 8'd135}: color_data = 12'hfff;
			{8'd97, 8'd136}: color_data = 12'hfff;
			{8'd97, 8'd137}: color_data = 12'hfff;
			{8'd97, 8'd138}: color_data = 12'hfff;
			{8'd97, 8'd139}: color_data = 12'haaa;
			{8'd97, 8'd140}: color_data = 12'h555;
			{8'd98, 8'd32}: color_data = 12'hd21;
			{8'd98, 8'd33}: color_data = 12'hd31;
			{8'd98, 8'd34}: color_data = 12'he31;
			{8'd98, 8'd35}: color_data = 12'he41;
			{8'd98, 8'd36}: color_data = 12'he41;
			{8'd98, 8'd37}: color_data = 12'he51;
			{8'd98, 8'd38}: color_data = 12'he51;
			{8'd98, 8'd39}: color_data = 12'he51;
			{8'd98, 8'd40}: color_data = 12'he61;
			{8'd98, 8'd41}: color_data = 12'he61;
			{8'd98, 8'd42}: color_data = 12'he71;
			{8'd98, 8'd43}: color_data = 12'he71;
			{8'd98, 8'd44}: color_data = 12'he71;
			{8'd98, 8'd45}: color_data = 12'he80;
			{8'd98, 8'd46}: color_data = 12'he80;
			{8'd98, 8'd47}: color_data = 12'he80;
			{8'd98, 8'd48}: color_data = 12'he90;
			{8'd98, 8'd49}: color_data = 12'he90;
			{8'd98, 8'd50}: color_data = 12'he90;
			{8'd98, 8'd51}: color_data = 12'hea0;
			{8'd98, 8'd52}: color_data = 12'hea0;
			{8'd98, 8'd53}: color_data = 12'h458;
			{8'd98, 8'd54}: color_data = 12'h677;
			{8'd98, 8'd55}: color_data = 12'h777;
			{8'd98, 8'd56}: color_data = 12'h666;
			{8'd98, 8'd57}: color_data = 12'h666;
			{8'd98, 8'd58}: color_data = 12'h666;
			{8'd98, 8'd59}: color_data = 12'h666;
			{8'd98, 8'd60}: color_data = 12'h666;
			{8'd98, 8'd61}: color_data = 12'h666;
			{8'd98, 8'd62}: color_data = 12'h666;
			{8'd98, 8'd63}: color_data = 12'h666;
			{8'd98, 8'd64}: color_data = 12'h666;
			{8'd98, 8'd65}: color_data = 12'h666;
			{8'd98, 8'd66}: color_data = 12'h666;
			{8'd98, 8'd67}: color_data = 12'h666;
			{8'd98, 8'd68}: color_data = 12'h555;
			{8'd98, 8'd69}: color_data = 12'h555;
			{8'd98, 8'd70}: color_data = 12'h555;
			{8'd98, 8'd71}: color_data = 12'h555;
			{8'd98, 8'd72}: color_data = 12'h555;
			{8'd98, 8'd73}: color_data = 12'h555;
			{8'd98, 8'd74}: color_data = 12'h555;
			{8'd98, 8'd75}: color_data = 12'h555;
			{8'd98, 8'd76}: color_data = 12'h555;
			{8'd98, 8'd77}: color_data = 12'h555;
			{8'd98, 8'd78}: color_data = 12'h555;
			{8'd98, 8'd79}: color_data = 12'h555;
			{8'd98, 8'd80}: color_data = 12'h555;
			{8'd98, 8'd81}: color_data = 12'h444;
			{8'd98, 8'd82}: color_data = 12'h444;
			{8'd98, 8'd83}: color_data = 12'h444;
			{8'd98, 8'd84}: color_data = 12'h444;
			{8'd98, 8'd85}: color_data = 12'h444;
			{8'd98, 8'd86}: color_data = 12'h444;
			{8'd98, 8'd87}: color_data = 12'h444;
			{8'd98, 8'd88}: color_data = 12'h444;
			{8'd98, 8'd89}: color_data = 12'h444;
			{8'd98, 8'd90}: color_data = 12'h444;
			{8'd98, 8'd91}: color_data = 12'h444;
			{8'd98, 8'd92}: color_data = 12'h444;
			{8'd98, 8'd93}: color_data = 12'h444;
			{8'd98, 8'd94}: color_data = 12'h333;
			{8'd98, 8'd95}: color_data = 12'h333;
			{8'd98, 8'd96}: color_data = 12'h333;
			{8'd98, 8'd97}: color_data = 12'h333;
			{8'd98, 8'd98}: color_data = 12'h333;
			{8'd98, 8'd99}: color_data = 12'h333;
			{8'd98, 8'd100}: color_data = 12'h333;
			{8'd98, 8'd101}: color_data = 12'h333;
			{8'd98, 8'd102}: color_data = 12'h333;
			{8'd98, 8'd103}: color_data = 12'h333;
			{8'd98, 8'd104}: color_data = 12'h333;
			{8'd98, 8'd105}: color_data = 12'h333;
			{8'd98, 8'd106}: color_data = 12'h333;
			{8'd98, 8'd107}: color_data = 12'h222;
			{8'd98, 8'd108}: color_data = 12'h222;
			{8'd98, 8'd109}: color_data = 12'h222;
			{8'd98, 8'd110}: color_data = 12'h222;
			{8'd98, 8'd111}: color_data = 12'h222;
			{8'd98, 8'd112}: color_data = 12'h222;
			{8'd98, 8'd113}: color_data = 12'h222;
			{8'd98, 8'd114}: color_data = 12'h222;
			{8'd98, 8'd115}: color_data = 12'h222;
			{8'd98, 8'd116}: color_data = 12'h222;
			{8'd98, 8'd117}: color_data = 12'h222;
			{8'd98, 8'd118}: color_data = 12'h222;
			{8'd98, 8'd119}: color_data = 12'h222;
			{8'd98, 8'd120}: color_data = 12'h222;
			{8'd98, 8'd121}: color_data = 12'h111;
			{8'd98, 8'd122}: color_data = 12'h111;
			{8'd98, 8'd123}: color_data = 12'h333;
			{8'd98, 8'd124}: color_data = 12'hccc;
			{8'd98, 8'd125}: color_data = 12'hfff;
			{8'd98, 8'd126}: color_data = 12'hfff;
			{8'd98, 8'd127}: color_data = 12'hfff;
			{8'd98, 8'd128}: color_data = 12'hfff;
			{8'd98, 8'd129}: color_data = 12'hfff;
			{8'd98, 8'd130}: color_data = 12'hfff;
			{8'd98, 8'd131}: color_data = 12'hfff;
			{8'd98, 8'd132}: color_data = 12'hfff;
			{8'd98, 8'd133}: color_data = 12'hfff;
			{8'd98, 8'd134}: color_data = 12'hfff;
			{8'd98, 8'd135}: color_data = 12'hfff;
			{8'd98, 8'd136}: color_data = 12'hfff;
			{8'd98, 8'd137}: color_data = 12'hfff;
			{8'd98, 8'd138}: color_data = 12'hfff;
			{8'd98, 8'd139}: color_data = 12'hbbb;
			{8'd98, 8'd140}: color_data = 12'h666;
			{8'd99, 8'd32}: color_data = 12'hb21;
			{8'd99, 8'd33}: color_data = 12'hc21;
			{8'd99, 8'd34}: color_data = 12'he31;
			{8'd99, 8'd35}: color_data = 12'he41;
			{8'd99, 8'd36}: color_data = 12'he41;
			{8'd99, 8'd37}: color_data = 12'he51;
			{8'd99, 8'd38}: color_data = 12'he51;
			{8'd99, 8'd39}: color_data = 12'he51;
			{8'd99, 8'd40}: color_data = 12'he61;
			{8'd99, 8'd41}: color_data = 12'he61;
			{8'd99, 8'd42}: color_data = 12'he71;
			{8'd99, 8'd43}: color_data = 12'he71;
			{8'd99, 8'd44}: color_data = 12'he71;
			{8'd99, 8'd45}: color_data = 12'hd70;
			{8'd99, 8'd46}: color_data = 12'hd80;
			{8'd99, 8'd47}: color_data = 12'he80;
			{8'd99, 8'd48}: color_data = 12'he90;
			{8'd99, 8'd49}: color_data = 12'he90;
			{8'd99, 8'd50}: color_data = 12'he90;
			{8'd99, 8'd51}: color_data = 12'he90;
			{8'd99, 8'd52}: color_data = 12'hea0;
			{8'd99, 8'd53}: color_data = 12'h667;
			{8'd99, 8'd54}: color_data = 12'h777;
			{8'd99, 8'd55}: color_data = 12'h777;
			{8'd99, 8'd56}: color_data = 12'h666;
			{8'd99, 8'd57}: color_data = 12'h666;
			{8'd99, 8'd58}: color_data = 12'h666;
			{8'd99, 8'd59}: color_data = 12'h666;
			{8'd99, 8'd60}: color_data = 12'h666;
			{8'd99, 8'd61}: color_data = 12'h666;
			{8'd99, 8'd62}: color_data = 12'h666;
			{8'd99, 8'd63}: color_data = 12'h666;
			{8'd99, 8'd64}: color_data = 12'h666;
			{8'd99, 8'd65}: color_data = 12'h666;
			{8'd99, 8'd66}: color_data = 12'h666;
			{8'd99, 8'd67}: color_data = 12'h666;
			{8'd99, 8'd68}: color_data = 12'h555;
			{8'd99, 8'd69}: color_data = 12'h555;
			{8'd99, 8'd70}: color_data = 12'h555;
			{8'd99, 8'd71}: color_data = 12'h555;
			{8'd99, 8'd72}: color_data = 12'h555;
			{8'd99, 8'd73}: color_data = 12'h555;
			{8'd99, 8'd74}: color_data = 12'h555;
			{8'd99, 8'd75}: color_data = 12'h555;
			{8'd99, 8'd76}: color_data = 12'h555;
			{8'd99, 8'd77}: color_data = 12'h555;
			{8'd99, 8'd78}: color_data = 12'h555;
			{8'd99, 8'd79}: color_data = 12'h555;
			{8'd99, 8'd80}: color_data = 12'h555;
			{8'd99, 8'd81}: color_data = 12'h444;
			{8'd99, 8'd82}: color_data = 12'h444;
			{8'd99, 8'd83}: color_data = 12'h444;
			{8'd99, 8'd84}: color_data = 12'h444;
			{8'd99, 8'd85}: color_data = 12'h444;
			{8'd99, 8'd86}: color_data = 12'h444;
			{8'd99, 8'd87}: color_data = 12'h444;
			{8'd99, 8'd88}: color_data = 12'h444;
			{8'd99, 8'd89}: color_data = 12'h444;
			{8'd99, 8'd90}: color_data = 12'h444;
			{8'd99, 8'd91}: color_data = 12'h444;
			{8'd99, 8'd92}: color_data = 12'h444;
			{8'd99, 8'd93}: color_data = 12'h444;
			{8'd99, 8'd94}: color_data = 12'h333;
			{8'd99, 8'd95}: color_data = 12'h333;
			{8'd99, 8'd96}: color_data = 12'h333;
			{8'd99, 8'd97}: color_data = 12'h333;
			{8'd99, 8'd98}: color_data = 12'h333;
			{8'd99, 8'd99}: color_data = 12'h333;
			{8'd99, 8'd100}: color_data = 12'h333;
			{8'd99, 8'd101}: color_data = 12'h333;
			{8'd99, 8'd102}: color_data = 12'h333;
			{8'd99, 8'd103}: color_data = 12'h333;
			{8'd99, 8'd104}: color_data = 12'h333;
			{8'd99, 8'd105}: color_data = 12'h333;
			{8'd99, 8'd106}: color_data = 12'h333;
			{8'd99, 8'd107}: color_data = 12'h222;
			{8'd99, 8'd108}: color_data = 12'h222;
			{8'd99, 8'd109}: color_data = 12'h222;
			{8'd99, 8'd110}: color_data = 12'h222;
			{8'd99, 8'd111}: color_data = 12'h222;
			{8'd99, 8'd112}: color_data = 12'h222;
			{8'd99, 8'd113}: color_data = 12'h222;
			{8'd99, 8'd114}: color_data = 12'h222;
			{8'd99, 8'd115}: color_data = 12'h222;
			{8'd99, 8'd116}: color_data = 12'h222;
			{8'd99, 8'd117}: color_data = 12'h222;
			{8'd99, 8'd118}: color_data = 12'h222;
			{8'd99, 8'd119}: color_data = 12'h222;
			{8'd99, 8'd120}: color_data = 12'h222;
			{8'd99, 8'd121}: color_data = 12'h111;
			{8'd99, 8'd122}: color_data = 12'h111;
			{8'd99, 8'd123}: color_data = 12'h444;
			{8'd99, 8'd124}: color_data = 12'hddd;
			{8'd99, 8'd125}: color_data = 12'hfff;
			{8'd99, 8'd126}: color_data = 12'hfff;
			{8'd99, 8'd127}: color_data = 12'hfff;
			{8'd99, 8'd128}: color_data = 12'hfff;
			{8'd99, 8'd129}: color_data = 12'hfff;
			{8'd99, 8'd130}: color_data = 12'hfff;
			{8'd99, 8'd131}: color_data = 12'hfff;
			{8'd99, 8'd132}: color_data = 12'hfff;
			{8'd99, 8'd133}: color_data = 12'hfff;
			{8'd99, 8'd134}: color_data = 12'hfff;
			{8'd99, 8'd135}: color_data = 12'hfff;
			{8'd99, 8'd136}: color_data = 12'hfff;
			{8'd99, 8'd137}: color_data = 12'hfff;
			{8'd99, 8'd138}: color_data = 12'hfff;
			{8'd99, 8'd139}: color_data = 12'hccc;
			{8'd99, 8'd140}: color_data = 12'h888;
			{8'd100, 8'd27}: color_data = 12'h777;
			{8'd100, 8'd28}: color_data = 12'h999;
			{8'd100, 8'd29}: color_data = 12'h888;
			{8'd100, 8'd30}: color_data = 12'h888;
			{8'd100, 8'd31}: color_data = 12'h789;
			{8'd100, 8'd32}: color_data = 12'hc20;
			{8'd100, 8'd33}: color_data = 12'hd31;
			{8'd100, 8'd34}: color_data = 12'hd31;
			{8'd100, 8'd35}: color_data = 12'he41;
			{8'd100, 8'd36}: color_data = 12'he41;
			{8'd100, 8'd37}: color_data = 12'hd51;
			{8'd100, 8'd38}: color_data = 12'hc51;
			{8'd100, 8'd39}: color_data = 12'hd51;
			{8'd100, 8'd40}: color_data = 12'he61;
			{8'd100, 8'd41}: color_data = 12'he61;
			{8'd100, 8'd42}: color_data = 12'he71;
			{8'd100, 8'd43}: color_data = 12'he71;
			{8'd100, 8'd44}: color_data = 12'hd71;
			{8'd100, 8'd45}: color_data = 12'hb60;
			{8'd100, 8'd46}: color_data = 12'hc70;
			{8'd100, 8'd47}: color_data = 12'he80;
			{8'd100, 8'd48}: color_data = 12'he90;
			{8'd100, 8'd49}: color_data = 12'he90;
			{8'd100, 8'd50}: color_data = 12'he90;
			{8'd100, 8'd51}: color_data = 12'hea0;
			{8'd100, 8'd52}: color_data = 12'hea0;
			{8'd100, 8'd53}: color_data = 12'h667;
			{8'd100, 8'd54}: color_data = 12'h777;
			{8'd100, 8'd55}: color_data = 12'h777;
			{8'd100, 8'd56}: color_data = 12'h666;
			{8'd100, 8'd57}: color_data = 12'h666;
			{8'd100, 8'd58}: color_data = 12'h666;
			{8'd100, 8'd59}: color_data = 12'h666;
			{8'd100, 8'd60}: color_data = 12'h666;
			{8'd100, 8'd61}: color_data = 12'h666;
			{8'd100, 8'd62}: color_data = 12'h666;
			{8'd100, 8'd63}: color_data = 12'h666;
			{8'd100, 8'd64}: color_data = 12'h666;
			{8'd100, 8'd65}: color_data = 12'h666;
			{8'd100, 8'd66}: color_data = 12'h666;
			{8'd100, 8'd67}: color_data = 12'h666;
			{8'd100, 8'd68}: color_data = 12'h555;
			{8'd100, 8'd69}: color_data = 12'h555;
			{8'd100, 8'd70}: color_data = 12'h555;
			{8'd100, 8'd71}: color_data = 12'h555;
			{8'd100, 8'd72}: color_data = 12'h555;
			{8'd100, 8'd73}: color_data = 12'h555;
			{8'd100, 8'd74}: color_data = 12'h555;
			{8'd100, 8'd75}: color_data = 12'h555;
			{8'd100, 8'd76}: color_data = 12'h555;
			{8'd100, 8'd77}: color_data = 12'h555;
			{8'd100, 8'd78}: color_data = 12'h555;
			{8'd100, 8'd79}: color_data = 12'h555;
			{8'd100, 8'd80}: color_data = 12'h555;
			{8'd100, 8'd81}: color_data = 12'h444;
			{8'd100, 8'd82}: color_data = 12'h444;
			{8'd100, 8'd83}: color_data = 12'h444;
			{8'd100, 8'd84}: color_data = 12'h444;
			{8'd100, 8'd85}: color_data = 12'h444;
			{8'd100, 8'd86}: color_data = 12'h444;
			{8'd100, 8'd87}: color_data = 12'h444;
			{8'd100, 8'd88}: color_data = 12'h444;
			{8'd100, 8'd89}: color_data = 12'h444;
			{8'd100, 8'd90}: color_data = 12'h444;
			{8'd100, 8'd91}: color_data = 12'h444;
			{8'd100, 8'd92}: color_data = 12'h444;
			{8'd100, 8'd93}: color_data = 12'h444;
			{8'd100, 8'd94}: color_data = 12'h333;
			{8'd100, 8'd95}: color_data = 12'h333;
			{8'd100, 8'd96}: color_data = 12'h333;
			{8'd100, 8'd97}: color_data = 12'h333;
			{8'd100, 8'd98}: color_data = 12'h333;
			{8'd100, 8'd99}: color_data = 12'h333;
			{8'd100, 8'd100}: color_data = 12'h333;
			{8'd100, 8'd101}: color_data = 12'h333;
			{8'd100, 8'd102}: color_data = 12'h333;
			{8'd100, 8'd103}: color_data = 12'h333;
			{8'd100, 8'd104}: color_data = 12'h333;
			{8'd100, 8'd105}: color_data = 12'h333;
			{8'd100, 8'd106}: color_data = 12'h333;
			{8'd100, 8'd107}: color_data = 12'h222;
			{8'd100, 8'd108}: color_data = 12'h222;
			{8'd100, 8'd109}: color_data = 12'h222;
			{8'd100, 8'd110}: color_data = 12'h222;
			{8'd100, 8'd111}: color_data = 12'h222;
			{8'd100, 8'd112}: color_data = 12'h222;
			{8'd100, 8'd113}: color_data = 12'h222;
			{8'd100, 8'd114}: color_data = 12'h222;
			{8'd100, 8'd115}: color_data = 12'h222;
			{8'd100, 8'd116}: color_data = 12'h222;
			{8'd100, 8'd117}: color_data = 12'h222;
			{8'd100, 8'd118}: color_data = 12'h222;
			{8'd100, 8'd119}: color_data = 12'h222;
			{8'd100, 8'd120}: color_data = 12'h222;
			{8'd100, 8'd121}: color_data = 12'h111;
			{8'd100, 8'd122}: color_data = 12'h111;
			{8'd100, 8'd123}: color_data = 12'h555;
			{8'd100, 8'd124}: color_data = 12'heee;
			{8'd100, 8'd125}: color_data = 12'hfff;
			{8'd100, 8'd126}: color_data = 12'hfff;
			{8'd100, 8'd127}: color_data = 12'hfff;
			{8'd100, 8'd128}: color_data = 12'hfff;
			{8'd100, 8'd129}: color_data = 12'hfff;
			{8'd100, 8'd130}: color_data = 12'hfff;
			{8'd100, 8'd131}: color_data = 12'hfff;
			{8'd100, 8'd132}: color_data = 12'hfff;
			{8'd100, 8'd133}: color_data = 12'hfff;
			{8'd100, 8'd134}: color_data = 12'hfff;
			{8'd100, 8'd135}: color_data = 12'hfff;
			{8'd100, 8'd136}: color_data = 12'hfff;
			{8'd100, 8'd137}: color_data = 12'hfff;
			{8'd100, 8'd138}: color_data = 12'hfff;
			{8'd100, 8'd139}: color_data = 12'hddd;
			{8'd100, 8'd140}: color_data = 12'haaa;
			{8'd101, 8'd22}: color_data = 12'h999;
			{8'd101, 8'd23}: color_data = 12'h988;
			{8'd101, 8'd24}: color_data = 12'h999;
			{8'd101, 8'd25}: color_data = 12'h999;
			{8'd101, 8'd26}: color_data = 12'h999;
			{8'd101, 8'd27}: color_data = 12'h999;
			{8'd101, 8'd28}: color_data = 12'h999;
			{8'd101, 8'd29}: color_data = 12'h999;
			{8'd101, 8'd30}: color_data = 12'h888;
			{8'd101, 8'd31}: color_data = 12'h788;
			{8'd101, 8'd32}: color_data = 12'hc20;
			{8'd101, 8'd33}: color_data = 12'hd31;
			{8'd101, 8'd34}: color_data = 12'hd31;
			{8'd101, 8'd35}: color_data = 12'hd41;
			{8'd101, 8'd36}: color_data = 12'he41;
			{8'd101, 8'd37}: color_data = 12'hc41;
			{8'd101, 8'd38}: color_data = 12'h830;
			{8'd101, 8'd39}: color_data = 12'hb40;
			{8'd101, 8'd40}: color_data = 12'he61;
			{8'd101, 8'd41}: color_data = 12'he61;
			{8'd101, 8'd42}: color_data = 12'he71;
			{8'd101, 8'd43}: color_data = 12'he71;
			{8'd101, 8'd44}: color_data = 12'he71;
			{8'd101, 8'd46}: color_data = 12'hc70;
			{8'd101, 8'd47}: color_data = 12'he80;
			{8'd101, 8'd48}: color_data = 12'he90;
			{8'd101, 8'd49}: color_data = 12'he90;
			{8'd101, 8'd50}: color_data = 12'he90;
			{8'd101, 8'd51}: color_data = 12'he90;
			{8'd101, 8'd52}: color_data = 12'he90;
			{8'd101, 8'd53}: color_data = 12'h667;
			{8'd101, 8'd54}: color_data = 12'h777;
			{8'd101, 8'd55}: color_data = 12'h777;
			{8'd101, 8'd56}: color_data = 12'h666;
			{8'd101, 8'd57}: color_data = 12'h666;
			{8'd101, 8'd58}: color_data = 12'h666;
			{8'd101, 8'd59}: color_data = 12'h666;
			{8'd101, 8'd60}: color_data = 12'h666;
			{8'd101, 8'd61}: color_data = 12'h666;
			{8'd101, 8'd62}: color_data = 12'h666;
			{8'd101, 8'd63}: color_data = 12'h666;
			{8'd101, 8'd64}: color_data = 12'h666;
			{8'd101, 8'd65}: color_data = 12'h666;
			{8'd101, 8'd66}: color_data = 12'h666;
			{8'd101, 8'd67}: color_data = 12'h666;
			{8'd101, 8'd68}: color_data = 12'h666;
			{8'd101, 8'd69}: color_data = 12'h555;
			{8'd101, 8'd70}: color_data = 12'h555;
			{8'd101, 8'd71}: color_data = 12'h555;
			{8'd101, 8'd72}: color_data = 12'h555;
			{8'd101, 8'd73}: color_data = 12'h555;
			{8'd101, 8'd74}: color_data = 12'h555;
			{8'd101, 8'd75}: color_data = 12'h555;
			{8'd101, 8'd76}: color_data = 12'h555;
			{8'd101, 8'd77}: color_data = 12'h555;
			{8'd101, 8'd78}: color_data = 12'h555;
			{8'd101, 8'd79}: color_data = 12'h555;
			{8'd101, 8'd80}: color_data = 12'h555;
			{8'd101, 8'd81}: color_data = 12'h444;
			{8'd101, 8'd82}: color_data = 12'h444;
			{8'd101, 8'd83}: color_data = 12'h444;
			{8'd101, 8'd84}: color_data = 12'h444;
			{8'd101, 8'd85}: color_data = 12'h444;
			{8'd101, 8'd86}: color_data = 12'h444;
			{8'd101, 8'd87}: color_data = 12'h444;
			{8'd101, 8'd88}: color_data = 12'h444;
			{8'd101, 8'd89}: color_data = 12'h444;
			{8'd101, 8'd90}: color_data = 12'h444;
			{8'd101, 8'd91}: color_data = 12'h444;
			{8'd101, 8'd92}: color_data = 12'h444;
			{8'd101, 8'd93}: color_data = 12'h444;
			{8'd101, 8'd94}: color_data = 12'h333;
			{8'd101, 8'd95}: color_data = 12'h333;
			{8'd101, 8'd96}: color_data = 12'h333;
			{8'd101, 8'd97}: color_data = 12'h333;
			{8'd101, 8'd98}: color_data = 12'h333;
			{8'd101, 8'd99}: color_data = 12'h333;
			{8'd101, 8'd100}: color_data = 12'h333;
			{8'd101, 8'd101}: color_data = 12'h333;
			{8'd101, 8'd102}: color_data = 12'h333;
			{8'd101, 8'd103}: color_data = 12'h333;
			{8'd101, 8'd104}: color_data = 12'h333;
			{8'd101, 8'd105}: color_data = 12'h333;
			{8'd101, 8'd106}: color_data = 12'h333;
			{8'd101, 8'd107}: color_data = 12'h222;
			{8'd101, 8'd108}: color_data = 12'h222;
			{8'd101, 8'd109}: color_data = 12'h222;
			{8'd101, 8'd110}: color_data = 12'h222;
			{8'd101, 8'd111}: color_data = 12'h222;
			{8'd101, 8'd112}: color_data = 12'h222;
			{8'd101, 8'd113}: color_data = 12'h222;
			{8'd101, 8'd114}: color_data = 12'h222;
			{8'd101, 8'd115}: color_data = 12'h222;
			{8'd101, 8'd116}: color_data = 12'h222;
			{8'd101, 8'd117}: color_data = 12'h222;
			{8'd101, 8'd118}: color_data = 12'h222;
			{8'd101, 8'd119}: color_data = 12'h222;
			{8'd101, 8'd120}: color_data = 12'h222;
			{8'd101, 8'd121}: color_data = 12'h111;
			{8'd101, 8'd122}: color_data = 12'h111;
			{8'd101, 8'd123}: color_data = 12'h666;
			{8'd101, 8'd124}: color_data = 12'hfff;
			{8'd101, 8'd125}: color_data = 12'hfff;
			{8'd101, 8'd126}: color_data = 12'hfff;
			{8'd101, 8'd127}: color_data = 12'hfff;
			{8'd101, 8'd128}: color_data = 12'hfff;
			{8'd101, 8'd129}: color_data = 12'hfff;
			{8'd101, 8'd130}: color_data = 12'hfff;
			{8'd101, 8'd131}: color_data = 12'hfff;
			{8'd101, 8'd132}: color_data = 12'hfff;
			{8'd101, 8'd133}: color_data = 12'hfff;
			{8'd101, 8'd134}: color_data = 12'hfff;
			{8'd101, 8'd135}: color_data = 12'hfff;
			{8'd101, 8'd136}: color_data = 12'hfff;
			{8'd101, 8'd137}: color_data = 12'hfff;
			{8'd101, 8'd138}: color_data = 12'hfff;
			{8'd101, 8'd139}: color_data = 12'heee;
			{8'd101, 8'd140}: color_data = 12'hbbb;
			{8'd102, 8'd16}: color_data = 12'h999;
			{8'd102, 8'd17}: color_data = 12'h999;
			{8'd102, 8'd18}: color_data = 12'haaa;
			{8'd102, 8'd19}: color_data = 12'h999;
			{8'd102, 8'd20}: color_data = 12'h999;
			{8'd102, 8'd21}: color_data = 12'h999;
			{8'd102, 8'd22}: color_data = 12'h999;
			{8'd102, 8'd23}: color_data = 12'h999;
			{8'd102, 8'd24}: color_data = 12'h999;
			{8'd102, 8'd25}: color_data = 12'h999;
			{8'd102, 8'd26}: color_data = 12'h999;
			{8'd102, 8'd27}: color_data = 12'h999;
			{8'd102, 8'd28}: color_data = 12'h999;
			{8'd102, 8'd29}: color_data = 12'h999;
			{8'd102, 8'd30}: color_data = 12'h888;
			{8'd102, 8'd31}: color_data = 12'h0ff;
			{8'd102, 8'd32}: color_data = 12'hc21;
			{8'd102, 8'd33}: color_data = 12'hd31;
			{8'd102, 8'd34}: color_data = 12'hd31;
			{8'd102, 8'd35}: color_data = 12'hd41;
			{8'd102, 8'd36}: color_data = 12'he41;
			{8'd102, 8'd37}: color_data = 12'hd41;
			{8'd102, 8'd38}: color_data = 12'h711;
			{8'd102, 8'd39}: color_data = 12'hc50;
			{8'd102, 8'd40}: color_data = 12'he61;
			{8'd102, 8'd41}: color_data = 12'he61;
			{8'd102, 8'd42}: color_data = 12'he71;
			{8'd102, 8'd43}: color_data = 12'he71;
			{8'd102, 8'd44}: color_data = 12'hd70;
			{8'd102, 8'd46}: color_data = 12'hd70;
			{8'd102, 8'd47}: color_data = 12'he80;
			{8'd102, 8'd48}: color_data = 12'he90;
			{8'd102, 8'd49}: color_data = 12'he90;
			{8'd102, 8'd50}: color_data = 12'he90;
			{8'd102, 8'd51}: color_data = 12'he90;
			{8'd102, 8'd52}: color_data = 12'he90;
			{8'd102, 8'd53}: color_data = 12'h677;
			{8'd102, 8'd54}: color_data = 12'h777;
			{8'd102, 8'd55}: color_data = 12'h777;
			{8'd102, 8'd56}: color_data = 12'h666;
			{8'd102, 8'd57}: color_data = 12'h666;
			{8'd102, 8'd58}: color_data = 12'h666;
			{8'd102, 8'd59}: color_data = 12'h666;
			{8'd102, 8'd60}: color_data = 12'h666;
			{8'd102, 8'd61}: color_data = 12'h666;
			{8'd102, 8'd62}: color_data = 12'h666;
			{8'd102, 8'd63}: color_data = 12'h666;
			{8'd102, 8'd64}: color_data = 12'h666;
			{8'd102, 8'd65}: color_data = 12'h666;
			{8'd102, 8'd66}: color_data = 12'h666;
			{8'd102, 8'd67}: color_data = 12'h666;
			{8'd102, 8'd68}: color_data = 12'h666;
			{8'd102, 8'd69}: color_data = 12'h555;
			{8'd102, 8'd70}: color_data = 12'h555;
			{8'd102, 8'd71}: color_data = 12'h555;
			{8'd102, 8'd72}: color_data = 12'h555;
			{8'd102, 8'd73}: color_data = 12'h555;
			{8'd102, 8'd74}: color_data = 12'h555;
			{8'd102, 8'd75}: color_data = 12'h555;
			{8'd102, 8'd76}: color_data = 12'h555;
			{8'd102, 8'd77}: color_data = 12'h555;
			{8'd102, 8'd78}: color_data = 12'h555;
			{8'd102, 8'd79}: color_data = 12'h555;
			{8'd102, 8'd80}: color_data = 12'h555;
			{8'd102, 8'd81}: color_data = 12'h444;
			{8'd102, 8'd82}: color_data = 12'h444;
			{8'd102, 8'd83}: color_data = 12'h444;
			{8'd102, 8'd84}: color_data = 12'h444;
			{8'd102, 8'd85}: color_data = 12'h444;
			{8'd102, 8'd86}: color_data = 12'h444;
			{8'd102, 8'd87}: color_data = 12'h444;
			{8'd102, 8'd88}: color_data = 12'h444;
			{8'd102, 8'd89}: color_data = 12'h444;
			{8'd102, 8'd90}: color_data = 12'h444;
			{8'd102, 8'd91}: color_data = 12'h444;
			{8'd102, 8'd92}: color_data = 12'h444;
			{8'd102, 8'd93}: color_data = 12'h444;
			{8'd102, 8'd94}: color_data = 12'h333;
			{8'd102, 8'd95}: color_data = 12'h333;
			{8'd102, 8'd96}: color_data = 12'h333;
			{8'd102, 8'd97}: color_data = 12'h333;
			{8'd102, 8'd98}: color_data = 12'h333;
			{8'd102, 8'd99}: color_data = 12'h333;
			{8'd102, 8'd100}: color_data = 12'h333;
			{8'd102, 8'd101}: color_data = 12'h333;
			{8'd102, 8'd102}: color_data = 12'h333;
			{8'd102, 8'd103}: color_data = 12'h333;
			{8'd102, 8'd104}: color_data = 12'h333;
			{8'd102, 8'd105}: color_data = 12'h333;
			{8'd102, 8'd106}: color_data = 12'h333;
			{8'd102, 8'd107}: color_data = 12'h333;
			{8'd102, 8'd108}: color_data = 12'h222;
			{8'd102, 8'd109}: color_data = 12'h222;
			{8'd102, 8'd110}: color_data = 12'h222;
			{8'd102, 8'd111}: color_data = 12'h222;
			{8'd102, 8'd112}: color_data = 12'h222;
			{8'd102, 8'd113}: color_data = 12'h222;
			{8'd102, 8'd114}: color_data = 12'h222;
			{8'd102, 8'd115}: color_data = 12'h222;
			{8'd102, 8'd116}: color_data = 12'h222;
			{8'd102, 8'd117}: color_data = 12'h222;
			{8'd102, 8'd118}: color_data = 12'h222;
			{8'd102, 8'd119}: color_data = 12'h222;
			{8'd102, 8'd120}: color_data = 12'h222;
			{8'd102, 8'd121}: color_data = 12'h111;
			{8'd102, 8'd122}: color_data = 12'h111;
			{8'd102, 8'd123}: color_data = 12'h888;
			{8'd102, 8'd124}: color_data = 12'hfff;
			{8'd102, 8'd125}: color_data = 12'hfff;
			{8'd102, 8'd126}: color_data = 12'hfff;
			{8'd102, 8'd127}: color_data = 12'hfff;
			{8'd102, 8'd128}: color_data = 12'hfff;
			{8'd102, 8'd129}: color_data = 12'hfff;
			{8'd102, 8'd130}: color_data = 12'hfff;
			{8'd102, 8'd131}: color_data = 12'hfff;
			{8'd102, 8'd132}: color_data = 12'hfff;
			{8'd102, 8'd133}: color_data = 12'hfff;
			{8'd102, 8'd134}: color_data = 12'hfff;
			{8'd102, 8'd135}: color_data = 12'hfff;
			{8'd102, 8'd136}: color_data = 12'hfff;
			{8'd102, 8'd137}: color_data = 12'hfff;
			{8'd102, 8'd138}: color_data = 12'hfff;
			{8'd102, 8'd139}: color_data = 12'heee;
			{8'd102, 8'd140}: color_data = 12'h999;
			{8'd102, 8'd141}: color_data = 12'h000;
			{8'd103, 8'd12}: color_data = 12'h999;
			{8'd103, 8'd13}: color_data = 12'h999;
			{8'd103, 8'd14}: color_data = 12'haaa;
			{8'd103, 8'd15}: color_data = 12'ha99;
			{8'd103, 8'd16}: color_data = 12'h999;
			{8'd103, 8'd17}: color_data = 12'h999;
			{8'd103, 8'd18}: color_data = 12'h999;
			{8'd103, 8'd19}: color_data = 12'h999;
			{8'd103, 8'd20}: color_data = 12'h999;
			{8'd103, 8'd21}: color_data = 12'h999;
			{8'd103, 8'd22}: color_data = 12'h999;
			{8'd103, 8'd23}: color_data = 12'h999;
			{8'd103, 8'd24}: color_data = 12'h999;
			{8'd103, 8'd25}: color_data = 12'h999;
			{8'd103, 8'd26}: color_data = 12'h999;
			{8'd103, 8'd27}: color_data = 12'h999;
			{8'd103, 8'd28}: color_data = 12'h999;
			{8'd103, 8'd29}: color_data = 12'h999;
			{8'd103, 8'd30}: color_data = 12'h888;
			{8'd103, 8'd32}: color_data = 12'hc21;
			{8'd103, 8'd33}: color_data = 12'he31;
			{8'd103, 8'd34}: color_data = 12'hd31;
			{8'd103, 8'd35}: color_data = 12'hd41;
			{8'd103, 8'd36}: color_data = 12'he41;
			{8'd103, 8'd37}: color_data = 12'hd41;
			{8'd103, 8'd38}: color_data = 12'hc31;
			{8'd103, 8'd39}: color_data = 12'hd61;
			{8'd103, 8'd40}: color_data = 12'he61;
			{8'd103, 8'd41}: color_data = 12'he61;
			{8'd103, 8'd42}: color_data = 12'he71;
			{8'd103, 8'd43}: color_data = 12'he71;
			{8'd103, 8'd44}: color_data = 12'hd70;
			{8'd103, 8'd45}: color_data = 12'hb30;
			{8'd103, 8'd46}: color_data = 12'hc70;
			{8'd103, 8'd47}: color_data = 12'he80;
			{8'd103, 8'd48}: color_data = 12'he90;
			{8'd103, 8'd49}: color_data = 12'he90;
			{8'd103, 8'd50}: color_data = 12'he90;
			{8'd103, 8'd51}: color_data = 12'hd90;
			{8'd103, 8'd52}: color_data = 12'hd90;
			{8'd103, 8'd53}: color_data = 12'h677;
			{8'd103, 8'd54}: color_data = 12'h777;
			{8'd103, 8'd55}: color_data = 12'h777;
			{8'd103, 8'd56}: color_data = 12'h666;
			{8'd103, 8'd57}: color_data = 12'h666;
			{8'd103, 8'd58}: color_data = 12'h666;
			{8'd103, 8'd59}: color_data = 12'h666;
			{8'd103, 8'd60}: color_data = 12'h666;
			{8'd103, 8'd61}: color_data = 12'h666;
			{8'd103, 8'd62}: color_data = 12'h666;
			{8'd103, 8'd63}: color_data = 12'h666;
			{8'd103, 8'd64}: color_data = 12'h666;
			{8'd103, 8'd65}: color_data = 12'h666;
			{8'd103, 8'd66}: color_data = 12'h666;
			{8'd103, 8'd67}: color_data = 12'h666;
			{8'd103, 8'd68}: color_data = 12'h666;
			{8'd103, 8'd69}: color_data = 12'h555;
			{8'd103, 8'd70}: color_data = 12'h555;
			{8'd103, 8'd71}: color_data = 12'h555;
			{8'd103, 8'd72}: color_data = 12'h555;
			{8'd103, 8'd73}: color_data = 12'h555;
			{8'd103, 8'd74}: color_data = 12'h555;
			{8'd103, 8'd75}: color_data = 12'h555;
			{8'd103, 8'd76}: color_data = 12'h555;
			{8'd103, 8'd77}: color_data = 12'h555;
			{8'd103, 8'd78}: color_data = 12'h555;
			{8'd103, 8'd79}: color_data = 12'h555;
			{8'd103, 8'd80}: color_data = 12'h555;
			{8'd103, 8'd81}: color_data = 12'h555;
			{8'd103, 8'd82}: color_data = 12'h444;
			{8'd103, 8'd83}: color_data = 12'h444;
			{8'd103, 8'd84}: color_data = 12'h444;
			{8'd103, 8'd85}: color_data = 12'h444;
			{8'd103, 8'd86}: color_data = 12'h444;
			{8'd103, 8'd87}: color_data = 12'h444;
			{8'd103, 8'd88}: color_data = 12'h444;
			{8'd103, 8'd89}: color_data = 12'h444;
			{8'd103, 8'd90}: color_data = 12'h444;
			{8'd103, 8'd91}: color_data = 12'h444;
			{8'd103, 8'd92}: color_data = 12'h444;
			{8'd103, 8'd93}: color_data = 12'h444;
			{8'd103, 8'd94}: color_data = 12'h444;
			{8'd103, 8'd95}: color_data = 12'h333;
			{8'd103, 8'd96}: color_data = 12'h333;
			{8'd103, 8'd97}: color_data = 12'h333;
			{8'd103, 8'd98}: color_data = 12'h333;
			{8'd103, 8'd99}: color_data = 12'h333;
			{8'd103, 8'd100}: color_data = 12'h333;
			{8'd103, 8'd101}: color_data = 12'h333;
			{8'd103, 8'd102}: color_data = 12'h333;
			{8'd103, 8'd103}: color_data = 12'h333;
			{8'd103, 8'd104}: color_data = 12'h333;
			{8'd103, 8'd105}: color_data = 12'h333;
			{8'd103, 8'd106}: color_data = 12'h333;
			{8'd103, 8'd107}: color_data = 12'h333;
			{8'd103, 8'd108}: color_data = 12'h222;
			{8'd103, 8'd109}: color_data = 12'h222;
			{8'd103, 8'd110}: color_data = 12'h222;
			{8'd103, 8'd111}: color_data = 12'h222;
			{8'd103, 8'd112}: color_data = 12'h222;
			{8'd103, 8'd113}: color_data = 12'h222;
			{8'd103, 8'd114}: color_data = 12'h222;
			{8'd103, 8'd115}: color_data = 12'h222;
			{8'd103, 8'd116}: color_data = 12'h222;
			{8'd103, 8'd117}: color_data = 12'h222;
			{8'd103, 8'd118}: color_data = 12'h222;
			{8'd103, 8'd119}: color_data = 12'h222;
			{8'd103, 8'd120}: color_data = 12'h222;
			{8'd103, 8'd121}: color_data = 12'h111;
			{8'd103, 8'd122}: color_data = 12'h222;
			{8'd103, 8'd123}: color_data = 12'h999;
			{8'd103, 8'd124}: color_data = 12'hfff;
			{8'd103, 8'd125}: color_data = 12'hfff;
			{8'd103, 8'd126}: color_data = 12'hfff;
			{8'd103, 8'd127}: color_data = 12'hfff;
			{8'd103, 8'd128}: color_data = 12'hfff;
			{8'd103, 8'd129}: color_data = 12'hfff;
			{8'd103, 8'd130}: color_data = 12'hfff;
			{8'd103, 8'd131}: color_data = 12'hfff;
			{8'd103, 8'd132}: color_data = 12'hfff;
			{8'd103, 8'd133}: color_data = 12'hfff;
			{8'd103, 8'd134}: color_data = 12'hfff;
			{8'd103, 8'd135}: color_data = 12'hfff;
			{8'd103, 8'd136}: color_data = 12'hfff;
			{8'd103, 8'd137}: color_data = 12'hfff;
			{8'd103, 8'd138}: color_data = 12'hfff;
			{8'd103, 8'd139}: color_data = 12'hfff;
			{8'd103, 8'd140}: color_data = 12'h999;
			{8'd103, 8'd141}: color_data = 12'h444;
			{8'd104, 8'd5}: color_data = 12'h000;
			{8'd104, 8'd6}: color_data = 12'haaa;
			{8'd104, 8'd7}: color_data = 12'haaa;
			{8'd104, 8'd8}: color_data = 12'haaa;
			{8'd104, 8'd9}: color_data = 12'haaa;
			{8'd104, 8'd10}: color_data = 12'haaa;
			{8'd104, 8'd11}: color_data = 12'haaa;
			{8'd104, 8'd12}: color_data = 12'haaa;
			{8'd104, 8'd13}: color_data = 12'haaa;
			{8'd104, 8'd14}: color_data = 12'haaa;
			{8'd104, 8'd15}: color_data = 12'haaa;
			{8'd104, 8'd16}: color_data = 12'haaa;
			{8'd104, 8'd17}: color_data = 12'haaa;
			{8'd104, 8'd18}: color_data = 12'haaa;
			{8'd104, 8'd19}: color_data = 12'h999;
			{8'd104, 8'd20}: color_data = 12'h999;
			{8'd104, 8'd21}: color_data = 12'h999;
			{8'd104, 8'd22}: color_data = 12'h999;
			{8'd104, 8'd23}: color_data = 12'h999;
			{8'd104, 8'd24}: color_data = 12'h999;
			{8'd104, 8'd25}: color_data = 12'h999;
			{8'd104, 8'd26}: color_data = 12'h999;
			{8'd104, 8'd27}: color_data = 12'h999;
			{8'd104, 8'd28}: color_data = 12'h999;
			{8'd104, 8'd29}: color_data = 12'h999;
			{8'd104, 8'd30}: color_data = 12'h888;
			{8'd104, 8'd31}: color_data = 12'hd00;
			{8'd104, 8'd32}: color_data = 12'hd21;
			{8'd104, 8'd33}: color_data = 12'he31;
			{8'd104, 8'd34}: color_data = 12'hd31;
			{8'd104, 8'd35}: color_data = 12'hd41;
			{8'd104, 8'd36}: color_data = 12'he41;
			{8'd104, 8'd37}: color_data = 12'hd41;
			{8'd104, 8'd38}: color_data = 12'hc41;
			{8'd104, 8'd39}: color_data = 12'hd51;
			{8'd104, 8'd40}: color_data = 12'he61;
			{8'd104, 8'd41}: color_data = 12'he61;
			{8'd104, 8'd42}: color_data = 12'he71;
			{8'd104, 8'd43}: color_data = 12'he71;
			{8'd104, 8'd44}: color_data = 12'hd70;
			{8'd104, 8'd45}: color_data = 12'hc61;
			{8'd104, 8'd46}: color_data = 12'hc70;
			{8'd104, 8'd47}: color_data = 12'he80;
			{8'd104, 8'd48}: color_data = 12'he90;
			{8'd104, 8'd49}: color_data = 12'he90;
			{8'd104, 8'd50}: color_data = 12'he90;
			{8'd104, 8'd51}: color_data = 12'hd90;
			{8'd104, 8'd52}: color_data = 12'hd90;
			{8'd104, 8'd53}: color_data = 12'h677;
			{8'd104, 8'd54}: color_data = 12'h777;
			{8'd104, 8'd55}: color_data = 12'h777;
			{8'd104, 8'd56}: color_data = 12'h666;
			{8'd104, 8'd57}: color_data = 12'h666;
			{8'd104, 8'd58}: color_data = 12'h666;
			{8'd104, 8'd59}: color_data = 12'h666;
			{8'd104, 8'd60}: color_data = 12'h666;
			{8'd104, 8'd61}: color_data = 12'h666;
			{8'd104, 8'd62}: color_data = 12'h666;
			{8'd104, 8'd63}: color_data = 12'h666;
			{8'd104, 8'd64}: color_data = 12'h666;
			{8'd104, 8'd65}: color_data = 12'h666;
			{8'd104, 8'd66}: color_data = 12'h666;
			{8'd104, 8'd67}: color_data = 12'h666;
			{8'd104, 8'd68}: color_data = 12'h666;
			{8'd104, 8'd69}: color_data = 12'h555;
			{8'd104, 8'd70}: color_data = 12'h555;
			{8'd104, 8'd71}: color_data = 12'h555;
			{8'd104, 8'd72}: color_data = 12'h555;
			{8'd104, 8'd73}: color_data = 12'h555;
			{8'd104, 8'd74}: color_data = 12'h555;
			{8'd104, 8'd75}: color_data = 12'h555;
			{8'd104, 8'd76}: color_data = 12'h555;
			{8'd104, 8'd77}: color_data = 12'h555;
			{8'd104, 8'd78}: color_data = 12'h555;
			{8'd104, 8'd79}: color_data = 12'h555;
			{8'd104, 8'd80}: color_data = 12'h555;
			{8'd104, 8'd81}: color_data = 12'h555;
			{8'd104, 8'd82}: color_data = 12'h444;
			{8'd104, 8'd83}: color_data = 12'h444;
			{8'd104, 8'd84}: color_data = 12'h444;
			{8'd104, 8'd85}: color_data = 12'h444;
			{8'd104, 8'd86}: color_data = 12'h444;
			{8'd104, 8'd87}: color_data = 12'h444;
			{8'd104, 8'd88}: color_data = 12'h444;
			{8'd104, 8'd89}: color_data = 12'h444;
			{8'd104, 8'd90}: color_data = 12'h444;
			{8'd104, 8'd91}: color_data = 12'h444;
			{8'd104, 8'd92}: color_data = 12'h444;
			{8'd104, 8'd93}: color_data = 12'h444;
			{8'd104, 8'd94}: color_data = 12'h444;
			{8'd104, 8'd95}: color_data = 12'h333;
			{8'd104, 8'd96}: color_data = 12'h333;
			{8'd104, 8'd97}: color_data = 12'h333;
			{8'd104, 8'd98}: color_data = 12'h333;
			{8'd104, 8'd99}: color_data = 12'h333;
			{8'd104, 8'd100}: color_data = 12'h333;
			{8'd104, 8'd101}: color_data = 12'h333;
			{8'd104, 8'd102}: color_data = 12'h333;
			{8'd104, 8'd103}: color_data = 12'h333;
			{8'd104, 8'd104}: color_data = 12'h333;
			{8'd104, 8'd105}: color_data = 12'h333;
			{8'd104, 8'd106}: color_data = 12'h333;
			{8'd104, 8'd107}: color_data = 12'h333;
			{8'd104, 8'd108}: color_data = 12'h222;
			{8'd104, 8'd109}: color_data = 12'h222;
			{8'd104, 8'd110}: color_data = 12'h222;
			{8'd104, 8'd111}: color_data = 12'h222;
			{8'd104, 8'd112}: color_data = 12'h222;
			{8'd104, 8'd113}: color_data = 12'h222;
			{8'd104, 8'd114}: color_data = 12'h222;
			{8'd104, 8'd115}: color_data = 12'h222;
			{8'd104, 8'd116}: color_data = 12'h222;
			{8'd104, 8'd117}: color_data = 12'h222;
			{8'd104, 8'd118}: color_data = 12'h222;
			{8'd104, 8'd119}: color_data = 12'h222;
			{8'd104, 8'd120}: color_data = 12'h222;
			{8'd104, 8'd121}: color_data = 12'h111;
			{8'd104, 8'd122}: color_data = 12'h222;
			{8'd104, 8'd123}: color_data = 12'haaa;
			{8'd104, 8'd124}: color_data = 12'hfff;
			{8'd104, 8'd125}: color_data = 12'hfff;
			{8'd104, 8'd126}: color_data = 12'hfff;
			{8'd104, 8'd127}: color_data = 12'hfff;
			{8'd104, 8'd128}: color_data = 12'hfff;
			{8'd104, 8'd129}: color_data = 12'hfff;
			{8'd104, 8'd130}: color_data = 12'hfff;
			{8'd104, 8'd131}: color_data = 12'hfff;
			{8'd104, 8'd132}: color_data = 12'hfff;
			{8'd104, 8'd133}: color_data = 12'hfff;
			{8'd104, 8'd134}: color_data = 12'hfff;
			{8'd104, 8'd135}: color_data = 12'hfff;
			{8'd104, 8'd136}: color_data = 12'hfff;
			{8'd104, 8'd137}: color_data = 12'hfff;
			{8'd104, 8'd138}: color_data = 12'hfff;
			{8'd104, 8'd139}: color_data = 12'hfff;
			{8'd104, 8'd140}: color_data = 12'h999;
			{8'd104, 8'd141}: color_data = 12'h555;
			{8'd105, 8'd1}: color_data = 12'hbbb;
			{8'd105, 8'd2}: color_data = 12'haaa;
			{8'd105, 8'd3}: color_data = 12'hbbb;
			{8'd105, 8'd4}: color_data = 12'haaa;
			{8'd105, 8'd5}: color_data = 12'haaa;
			{8'd105, 8'd6}: color_data = 12'haaa;
			{8'd105, 8'd7}: color_data = 12'haaa;
			{8'd105, 8'd8}: color_data = 12'haaa;
			{8'd105, 8'd9}: color_data = 12'haaa;
			{8'd105, 8'd10}: color_data = 12'haaa;
			{8'd105, 8'd11}: color_data = 12'haaa;
			{8'd105, 8'd12}: color_data = 12'haaa;
			{8'd105, 8'd13}: color_data = 12'haaa;
			{8'd105, 8'd14}: color_data = 12'haaa;
			{8'd105, 8'd15}: color_data = 12'haaa;
			{8'd105, 8'd16}: color_data = 12'haaa;
			{8'd105, 8'd17}: color_data = 12'h999;
			{8'd105, 8'd18}: color_data = 12'h999;
			{8'd105, 8'd19}: color_data = 12'h999;
			{8'd105, 8'd20}: color_data = 12'h999;
			{8'd105, 8'd21}: color_data = 12'h999;
			{8'd105, 8'd22}: color_data = 12'h999;
			{8'd105, 8'd23}: color_data = 12'h999;
			{8'd105, 8'd24}: color_data = 12'h999;
			{8'd105, 8'd25}: color_data = 12'h999;
			{8'd105, 8'd26}: color_data = 12'h999;
			{8'd105, 8'd27}: color_data = 12'h999;
			{8'd105, 8'd28}: color_data = 12'h999;
			{8'd105, 8'd29}: color_data = 12'h999;
			{8'd105, 8'd30}: color_data = 12'h899;
			{8'd105, 8'd31}: color_data = 12'hc00;
			{8'd105, 8'd32}: color_data = 12'hd21;
			{8'd105, 8'd33}: color_data = 12'he31;
			{8'd105, 8'd34}: color_data = 12'hd31;
			{8'd105, 8'd35}: color_data = 12'hd41;
			{8'd105, 8'd36}: color_data = 12'he41;
			{8'd105, 8'd37}: color_data = 12'hd41;
			{8'd105, 8'd38}: color_data = 12'hc41;
			{8'd105, 8'd39}: color_data = 12'hd51;
			{8'd105, 8'd40}: color_data = 12'he61;
			{8'd105, 8'd41}: color_data = 12'he61;
			{8'd105, 8'd42}: color_data = 12'he71;
			{8'd105, 8'd43}: color_data = 12'he71;
			{8'd105, 8'd44}: color_data = 12'hc60;
			{8'd105, 8'd45}: color_data = 12'ha40;
			{8'd105, 8'd46}: color_data = 12'hc70;
			{8'd105, 8'd47}: color_data = 12'hd80;
			{8'd105, 8'd48}: color_data = 12'he90;
			{8'd105, 8'd49}: color_data = 12'he90;
			{8'd105, 8'd50}: color_data = 12'he90;
			{8'd105, 8'd51}: color_data = 12'hd90;
			{8'd105, 8'd52}: color_data = 12'hd90;
			{8'd105, 8'd53}: color_data = 12'h677;
			{8'd105, 8'd54}: color_data = 12'h777;
			{8'd105, 8'd55}: color_data = 12'h777;
			{8'd105, 8'd56}: color_data = 12'h666;
			{8'd105, 8'd57}: color_data = 12'h666;
			{8'd105, 8'd58}: color_data = 12'h666;
			{8'd105, 8'd59}: color_data = 12'h666;
			{8'd105, 8'd60}: color_data = 12'h666;
			{8'd105, 8'd61}: color_data = 12'h666;
			{8'd105, 8'd62}: color_data = 12'h666;
			{8'd105, 8'd63}: color_data = 12'h666;
			{8'd105, 8'd64}: color_data = 12'h666;
			{8'd105, 8'd65}: color_data = 12'h666;
			{8'd105, 8'd66}: color_data = 12'h666;
			{8'd105, 8'd67}: color_data = 12'h666;
			{8'd105, 8'd68}: color_data = 12'h666;
			{8'd105, 8'd69}: color_data = 12'h555;
			{8'd105, 8'd70}: color_data = 12'h555;
			{8'd105, 8'd71}: color_data = 12'h555;
			{8'd105, 8'd72}: color_data = 12'h555;
			{8'd105, 8'd73}: color_data = 12'h555;
			{8'd105, 8'd74}: color_data = 12'h555;
			{8'd105, 8'd75}: color_data = 12'h555;
			{8'd105, 8'd76}: color_data = 12'h555;
			{8'd105, 8'd77}: color_data = 12'h555;
			{8'd105, 8'd78}: color_data = 12'h555;
			{8'd105, 8'd79}: color_data = 12'h555;
			{8'd105, 8'd80}: color_data = 12'h555;
			{8'd105, 8'd81}: color_data = 12'h555;
			{8'd105, 8'd82}: color_data = 12'h444;
			{8'd105, 8'd83}: color_data = 12'h444;
			{8'd105, 8'd84}: color_data = 12'h444;
			{8'd105, 8'd85}: color_data = 12'h444;
			{8'd105, 8'd86}: color_data = 12'h444;
			{8'd105, 8'd87}: color_data = 12'h444;
			{8'd105, 8'd88}: color_data = 12'h444;
			{8'd105, 8'd89}: color_data = 12'h444;
			{8'd105, 8'd90}: color_data = 12'h444;
			{8'd105, 8'd91}: color_data = 12'h444;
			{8'd105, 8'd92}: color_data = 12'h444;
			{8'd105, 8'd93}: color_data = 12'h444;
			{8'd105, 8'd94}: color_data = 12'h444;
			{8'd105, 8'd95}: color_data = 12'h333;
			{8'd105, 8'd96}: color_data = 12'h333;
			{8'd105, 8'd97}: color_data = 12'h333;
			{8'd105, 8'd98}: color_data = 12'h333;
			{8'd105, 8'd99}: color_data = 12'h333;
			{8'd105, 8'd100}: color_data = 12'h333;
			{8'd105, 8'd101}: color_data = 12'h333;
			{8'd105, 8'd102}: color_data = 12'h333;
			{8'd105, 8'd103}: color_data = 12'h333;
			{8'd105, 8'd104}: color_data = 12'h333;
			{8'd105, 8'd105}: color_data = 12'h333;
			{8'd105, 8'd106}: color_data = 12'h333;
			{8'd105, 8'd107}: color_data = 12'h333;
			{8'd105, 8'd108}: color_data = 12'h222;
			{8'd105, 8'd109}: color_data = 12'h222;
			{8'd105, 8'd110}: color_data = 12'h222;
			{8'd105, 8'd111}: color_data = 12'h222;
			{8'd105, 8'd112}: color_data = 12'h222;
			{8'd105, 8'd113}: color_data = 12'h222;
			{8'd105, 8'd114}: color_data = 12'h222;
			{8'd105, 8'd115}: color_data = 12'h222;
			{8'd105, 8'd116}: color_data = 12'h222;
			{8'd105, 8'd117}: color_data = 12'h222;
			{8'd105, 8'd118}: color_data = 12'h222;
			{8'd105, 8'd119}: color_data = 12'h222;
			{8'd105, 8'd120}: color_data = 12'h222;
			{8'd105, 8'd121}: color_data = 12'h111;
			{8'd105, 8'd122}: color_data = 12'h222;
			{8'd105, 8'd123}: color_data = 12'hbbb;
			{8'd105, 8'd124}: color_data = 12'hfff;
			{8'd105, 8'd125}: color_data = 12'hfff;
			{8'd105, 8'd126}: color_data = 12'hfff;
			{8'd105, 8'd127}: color_data = 12'hddd;
			{8'd105, 8'd128}: color_data = 12'haaa;
			{8'd105, 8'd129}: color_data = 12'haaa;
			{8'd105, 8'd130}: color_data = 12'hbbb;
			{8'd105, 8'd131}: color_data = 12'hfff;
			{8'd105, 8'd132}: color_data = 12'hfff;
			{8'd105, 8'd133}: color_data = 12'hfff;
			{8'd105, 8'd134}: color_data = 12'hfff;
			{8'd105, 8'd135}: color_data = 12'hfff;
			{8'd105, 8'd136}: color_data = 12'hfff;
			{8'd105, 8'd137}: color_data = 12'hfff;
			{8'd105, 8'd138}: color_data = 12'hfff;
			{8'd105, 8'd139}: color_data = 12'hfff;
			{8'd105, 8'd140}: color_data = 12'haaa;
			{8'd105, 8'd141}: color_data = 12'h777;
			{8'd106, 8'd0}: color_data = 12'hbbb;
			{8'd106, 8'd1}: color_data = 12'hbbb;
			{8'd106, 8'd2}: color_data = 12'hbbb;
			{8'd106, 8'd3}: color_data = 12'hbbb;
			{8'd106, 8'd4}: color_data = 12'hbbb;
			{8'd106, 8'd5}: color_data = 12'haaa;
			{8'd106, 8'd6}: color_data = 12'hbbb;
			{8'd106, 8'd7}: color_data = 12'hbbb;
			{8'd106, 8'd8}: color_data = 12'haaa;
			{8'd106, 8'd9}: color_data = 12'haaa;
			{8'd106, 8'd10}: color_data = 12'haaa;
			{8'd106, 8'd11}: color_data = 12'haaa;
			{8'd106, 8'd12}: color_data = 12'haaa;
			{8'd106, 8'd13}: color_data = 12'haaa;
			{8'd106, 8'd14}: color_data = 12'haaa;
			{8'd106, 8'd15}: color_data = 12'haaa;
			{8'd106, 8'd16}: color_data = 12'haaa;
			{8'd106, 8'd17}: color_data = 12'h999;
			{8'd106, 8'd18}: color_data = 12'h999;
			{8'd106, 8'd19}: color_data = 12'h999;
			{8'd106, 8'd20}: color_data = 12'h999;
			{8'd106, 8'd21}: color_data = 12'h999;
			{8'd106, 8'd22}: color_data = 12'h999;
			{8'd106, 8'd23}: color_data = 12'h999;
			{8'd106, 8'd24}: color_data = 12'h999;
			{8'd106, 8'd25}: color_data = 12'h999;
			{8'd106, 8'd26}: color_data = 12'h999;
			{8'd106, 8'd27}: color_data = 12'h999;
			{8'd106, 8'd28}: color_data = 12'h999;
			{8'd106, 8'd29}: color_data = 12'h888;
			{8'd106, 8'd30}: color_data = 12'h899;
			{8'd106, 8'd31}: color_data = 12'hc20;
			{8'd106, 8'd32}: color_data = 12'hd21;
			{8'd106, 8'd33}: color_data = 12'hd31;
			{8'd106, 8'd34}: color_data = 12'hd31;
			{8'd106, 8'd35}: color_data = 12'hd41;
			{8'd106, 8'd36}: color_data = 12'he41;
			{8'd106, 8'd37}: color_data = 12'hd41;
			{8'd106, 8'd38}: color_data = 12'hc40;
			{8'd106, 8'd39}: color_data = 12'hc51;
			{8'd106, 8'd40}: color_data = 12'hd61;
			{8'd106, 8'd41}: color_data = 12'hd61;
			{8'd106, 8'd42}: color_data = 12'hd61;
			{8'd106, 8'd43}: color_data = 12'hc60;
			{8'd106, 8'd44}: color_data = 12'hb60;
			{8'd106, 8'd46}: color_data = 12'hd70;
			{8'd106, 8'd47}: color_data = 12'he80;
			{8'd106, 8'd48}: color_data = 12'he90;
			{8'd106, 8'd49}: color_data = 12'he90;
			{8'd106, 8'd50}: color_data = 12'he90;
			{8'd106, 8'd51}: color_data = 12'hd90;
			{8'd106, 8'd52}: color_data = 12'hd90;
			{8'd106, 8'd53}: color_data = 12'h677;
			{8'd106, 8'd54}: color_data = 12'h777;
			{8'd106, 8'd55}: color_data = 12'h777;
			{8'd106, 8'd56}: color_data = 12'h666;
			{8'd106, 8'd57}: color_data = 12'h666;
			{8'd106, 8'd58}: color_data = 12'h666;
			{8'd106, 8'd59}: color_data = 12'h666;
			{8'd106, 8'd60}: color_data = 12'h666;
			{8'd106, 8'd61}: color_data = 12'h666;
			{8'd106, 8'd62}: color_data = 12'h666;
			{8'd106, 8'd63}: color_data = 12'h666;
			{8'd106, 8'd64}: color_data = 12'h666;
			{8'd106, 8'd65}: color_data = 12'h666;
			{8'd106, 8'd66}: color_data = 12'h666;
			{8'd106, 8'd67}: color_data = 12'h666;
			{8'd106, 8'd68}: color_data = 12'h666;
			{8'd106, 8'd69}: color_data = 12'h555;
			{8'd106, 8'd70}: color_data = 12'h555;
			{8'd106, 8'd71}: color_data = 12'h555;
			{8'd106, 8'd72}: color_data = 12'h555;
			{8'd106, 8'd73}: color_data = 12'h555;
			{8'd106, 8'd74}: color_data = 12'h555;
			{8'd106, 8'd75}: color_data = 12'h555;
			{8'd106, 8'd76}: color_data = 12'h555;
			{8'd106, 8'd77}: color_data = 12'h555;
			{8'd106, 8'd78}: color_data = 12'h555;
			{8'd106, 8'd79}: color_data = 12'h555;
			{8'd106, 8'd80}: color_data = 12'h555;
			{8'd106, 8'd81}: color_data = 12'h555;
			{8'd106, 8'd82}: color_data = 12'h444;
			{8'd106, 8'd83}: color_data = 12'h444;
			{8'd106, 8'd84}: color_data = 12'h444;
			{8'd106, 8'd85}: color_data = 12'h444;
			{8'd106, 8'd86}: color_data = 12'h444;
			{8'd106, 8'd87}: color_data = 12'h444;
			{8'd106, 8'd88}: color_data = 12'h444;
			{8'd106, 8'd89}: color_data = 12'h444;
			{8'd106, 8'd90}: color_data = 12'h444;
			{8'd106, 8'd91}: color_data = 12'h444;
			{8'd106, 8'd92}: color_data = 12'h444;
			{8'd106, 8'd93}: color_data = 12'h444;
			{8'd106, 8'd94}: color_data = 12'h444;
			{8'd106, 8'd95}: color_data = 12'h333;
			{8'd106, 8'd96}: color_data = 12'h333;
			{8'd106, 8'd97}: color_data = 12'h333;
			{8'd106, 8'd98}: color_data = 12'h333;
			{8'd106, 8'd99}: color_data = 12'h333;
			{8'd106, 8'd100}: color_data = 12'h333;
			{8'd106, 8'd101}: color_data = 12'h333;
			{8'd106, 8'd102}: color_data = 12'h333;
			{8'd106, 8'd103}: color_data = 12'h333;
			{8'd106, 8'd104}: color_data = 12'h333;
			{8'd106, 8'd105}: color_data = 12'h333;
			{8'd106, 8'd106}: color_data = 12'h333;
			{8'd106, 8'd107}: color_data = 12'h333;
			{8'd106, 8'd108}: color_data = 12'h222;
			{8'd106, 8'd109}: color_data = 12'h222;
			{8'd106, 8'd110}: color_data = 12'h222;
			{8'd106, 8'd111}: color_data = 12'h222;
			{8'd106, 8'd112}: color_data = 12'h222;
			{8'd106, 8'd113}: color_data = 12'h222;
			{8'd106, 8'd114}: color_data = 12'h222;
			{8'd106, 8'd115}: color_data = 12'h222;
			{8'd106, 8'd116}: color_data = 12'h222;
			{8'd106, 8'd117}: color_data = 12'h222;
			{8'd106, 8'd118}: color_data = 12'h222;
			{8'd106, 8'd119}: color_data = 12'h222;
			{8'd106, 8'd120}: color_data = 12'h222;
			{8'd106, 8'd121}: color_data = 12'h111;
			{8'd106, 8'd122}: color_data = 12'h222;
			{8'd106, 8'd123}: color_data = 12'hbbb;
			{8'd106, 8'd124}: color_data = 12'hfff;
			{8'd106, 8'd125}: color_data = 12'hfff;
			{8'd106, 8'd126}: color_data = 12'hcbc;
			{8'd106, 8'd127}: color_data = 12'h444;
			{8'd106, 8'd128}: color_data = 12'h432;
			{8'd106, 8'd129}: color_data = 12'h321;
			{8'd106, 8'd130}: color_data = 12'h554;
			{8'd106, 8'd131}: color_data = 12'hfff;
			{8'd106, 8'd132}: color_data = 12'hfff;
			{8'd106, 8'd133}: color_data = 12'hfff;
			{8'd106, 8'd134}: color_data = 12'hfff;
			{8'd106, 8'd135}: color_data = 12'hfff;
			{8'd106, 8'd136}: color_data = 12'hfff;
			{8'd106, 8'd137}: color_data = 12'hfff;
			{8'd106, 8'd138}: color_data = 12'hfff;
			{8'd106, 8'd139}: color_data = 12'hfff;
			{8'd106, 8'd140}: color_data = 12'hbbb;
			{8'd106, 8'd141}: color_data = 12'h888;
			{8'd107, 8'd0}: color_data = 12'hbbb;
			{8'd107, 8'd1}: color_data = 12'hbbb;
			{8'd107, 8'd2}: color_data = 12'hbbb;
			{8'd107, 8'd3}: color_data = 12'hbbb;
			{8'd107, 8'd4}: color_data = 12'hbbb;
			{8'd107, 8'd5}: color_data = 12'haaa;
			{8'd107, 8'd6}: color_data = 12'haaa;
			{8'd107, 8'd7}: color_data = 12'haaa;
			{8'd107, 8'd8}: color_data = 12'haaa;
			{8'd107, 8'd9}: color_data = 12'haaa;
			{8'd107, 8'd10}: color_data = 12'haaa;
			{8'd107, 8'd11}: color_data = 12'haaa;
			{8'd107, 8'd12}: color_data = 12'haaa;
			{8'd107, 8'd13}: color_data = 12'haaa;
			{8'd107, 8'd14}: color_data = 12'haaa;
			{8'd107, 8'd15}: color_data = 12'haaa;
			{8'd107, 8'd16}: color_data = 12'haaa;
			{8'd107, 8'd17}: color_data = 12'h999;
			{8'd107, 8'd18}: color_data = 12'h999;
			{8'd107, 8'd19}: color_data = 12'h999;
			{8'd107, 8'd20}: color_data = 12'h999;
			{8'd107, 8'd21}: color_data = 12'h999;
			{8'd107, 8'd22}: color_data = 12'h999;
			{8'd107, 8'd23}: color_data = 12'h999;
			{8'd107, 8'd24}: color_data = 12'h999;
			{8'd107, 8'd25}: color_data = 12'h999;
			{8'd107, 8'd26}: color_data = 12'h999;
			{8'd107, 8'd27}: color_data = 12'h999;
			{8'd107, 8'd28}: color_data = 12'h999;
			{8'd107, 8'd29}: color_data = 12'h888;
			{8'd107, 8'd30}: color_data = 12'h7ab;
			{8'd107, 8'd31}: color_data = 12'hd10;
			{8'd107, 8'd32}: color_data = 12'hd21;
			{8'd107, 8'd33}: color_data = 12'hd31;
			{8'd107, 8'd34}: color_data = 12'hd31;
			{8'd107, 8'd35}: color_data = 12'hd41;
			{8'd107, 8'd36}: color_data = 12'he41;
			{8'd107, 8'd37}: color_data = 12'hd41;
			{8'd107, 8'd38}: color_data = 12'hd40;
			{8'd107, 8'd40}: color_data = 12'hf00;
			{8'd107, 8'd41}: color_data = 12'hf20;
			{8'd107, 8'd42}: color_data = 12'hf20;
			{8'd107, 8'd43}: color_data = 12'hc00;
			{8'd107, 8'd44}: color_data = 12'hf00;
			{8'd107, 8'd46}: color_data = 12'he80;
			{8'd107, 8'd47}: color_data = 12'he80;
			{8'd107, 8'd48}: color_data = 12'he90;
			{8'd107, 8'd49}: color_data = 12'he90;
			{8'd107, 8'd50}: color_data = 12'he90;
			{8'd107, 8'd51}: color_data = 12'hd90;
			{8'd107, 8'd52}: color_data = 12'hd90;
			{8'd107, 8'd53}: color_data = 12'h677;
			{8'd107, 8'd54}: color_data = 12'h777;
			{8'd107, 8'd55}: color_data = 12'h777;
			{8'd107, 8'd56}: color_data = 12'h666;
			{8'd107, 8'd57}: color_data = 12'h666;
			{8'd107, 8'd58}: color_data = 12'h666;
			{8'd107, 8'd59}: color_data = 12'h666;
			{8'd107, 8'd60}: color_data = 12'h666;
			{8'd107, 8'd61}: color_data = 12'h666;
			{8'd107, 8'd62}: color_data = 12'h666;
			{8'd107, 8'd63}: color_data = 12'h666;
			{8'd107, 8'd64}: color_data = 12'h666;
			{8'd107, 8'd65}: color_data = 12'h666;
			{8'd107, 8'd66}: color_data = 12'h666;
			{8'd107, 8'd67}: color_data = 12'h666;
			{8'd107, 8'd68}: color_data = 12'h666;
			{8'd107, 8'd69}: color_data = 12'h555;
			{8'd107, 8'd70}: color_data = 12'h555;
			{8'd107, 8'd71}: color_data = 12'h555;
			{8'd107, 8'd72}: color_data = 12'h555;
			{8'd107, 8'd73}: color_data = 12'h555;
			{8'd107, 8'd74}: color_data = 12'h555;
			{8'd107, 8'd75}: color_data = 12'h555;
			{8'd107, 8'd76}: color_data = 12'h555;
			{8'd107, 8'd77}: color_data = 12'h555;
			{8'd107, 8'd78}: color_data = 12'h555;
			{8'd107, 8'd79}: color_data = 12'h555;
			{8'd107, 8'd80}: color_data = 12'h555;
			{8'd107, 8'd81}: color_data = 12'h555;
			{8'd107, 8'd82}: color_data = 12'h444;
			{8'd107, 8'd83}: color_data = 12'h444;
			{8'd107, 8'd84}: color_data = 12'h444;
			{8'd107, 8'd85}: color_data = 12'h444;
			{8'd107, 8'd86}: color_data = 12'h444;
			{8'd107, 8'd87}: color_data = 12'h444;
			{8'd107, 8'd88}: color_data = 12'h444;
			{8'd107, 8'd89}: color_data = 12'h444;
			{8'd107, 8'd90}: color_data = 12'h444;
			{8'd107, 8'd91}: color_data = 12'h444;
			{8'd107, 8'd92}: color_data = 12'h444;
			{8'd107, 8'd93}: color_data = 12'h444;
			{8'd107, 8'd94}: color_data = 12'h444;
			{8'd107, 8'd95}: color_data = 12'h333;
			{8'd107, 8'd96}: color_data = 12'h333;
			{8'd107, 8'd97}: color_data = 12'h333;
			{8'd107, 8'd98}: color_data = 12'h333;
			{8'd107, 8'd99}: color_data = 12'h333;
			{8'd107, 8'd100}: color_data = 12'h333;
			{8'd107, 8'd101}: color_data = 12'h333;
			{8'd107, 8'd102}: color_data = 12'h333;
			{8'd107, 8'd103}: color_data = 12'h333;
			{8'd107, 8'd104}: color_data = 12'h333;
			{8'd107, 8'd105}: color_data = 12'h333;
			{8'd107, 8'd106}: color_data = 12'h333;
			{8'd107, 8'd107}: color_data = 12'h333;
			{8'd107, 8'd108}: color_data = 12'h222;
			{8'd107, 8'd109}: color_data = 12'h222;
			{8'd107, 8'd110}: color_data = 12'h222;
			{8'd107, 8'd111}: color_data = 12'h222;
			{8'd107, 8'd112}: color_data = 12'h222;
			{8'd107, 8'd113}: color_data = 12'h222;
			{8'd107, 8'd114}: color_data = 12'h222;
			{8'd107, 8'd115}: color_data = 12'h222;
			{8'd107, 8'd116}: color_data = 12'h222;
			{8'd107, 8'd117}: color_data = 12'h222;
			{8'd107, 8'd118}: color_data = 12'h222;
			{8'd107, 8'd119}: color_data = 12'h222;
			{8'd107, 8'd120}: color_data = 12'h222;
			{8'd107, 8'd121}: color_data = 12'h111;
			{8'd107, 8'd122}: color_data = 12'h333;
			{8'd107, 8'd123}: color_data = 12'hccc;
			{8'd107, 8'd124}: color_data = 12'hfff;
			{8'd107, 8'd125}: color_data = 12'hcbb;
			{8'd107, 8'd126}: color_data = 12'h333;
			{8'd107, 8'd127}: color_data = 12'h532;
			{8'd107, 8'd128}: color_data = 12'h742;
			{8'd107, 8'd129}: color_data = 12'h531;
			{8'd107, 8'd130}: color_data = 12'h655;
			{8'd107, 8'd131}: color_data = 12'hfff;
			{8'd107, 8'd132}: color_data = 12'hfff;
			{8'd107, 8'd133}: color_data = 12'hfff;
			{8'd107, 8'd134}: color_data = 12'hfff;
			{8'd107, 8'd135}: color_data = 12'hfff;
			{8'd107, 8'd136}: color_data = 12'hfff;
			{8'd107, 8'd137}: color_data = 12'hfff;
			{8'd107, 8'd138}: color_data = 12'hfff;
			{8'd107, 8'd139}: color_data = 12'hfff;
			{8'd107, 8'd140}: color_data = 12'hccc;
			{8'd107, 8'd141}: color_data = 12'hbbb;
			{8'd108, 8'd0}: color_data = 12'hbbb;
			{8'd108, 8'd1}: color_data = 12'hbbb;
			{8'd108, 8'd2}: color_data = 12'hbbb;
			{8'd108, 8'd3}: color_data = 12'hbbb;
			{8'd108, 8'd4}: color_data = 12'haaa;
			{8'd108, 8'd5}: color_data = 12'haaa;
			{8'd108, 8'd6}: color_data = 12'haaa;
			{8'd108, 8'd7}: color_data = 12'haaa;
			{8'd108, 8'd8}: color_data = 12'haaa;
			{8'd108, 8'd9}: color_data = 12'haaa;
			{8'd108, 8'd10}: color_data = 12'haaa;
			{8'd108, 8'd11}: color_data = 12'haaa;
			{8'd108, 8'd12}: color_data = 12'haaa;
			{8'd108, 8'd13}: color_data = 12'haaa;
			{8'd108, 8'd14}: color_data = 12'haaa;
			{8'd108, 8'd15}: color_data = 12'haaa;
			{8'd108, 8'd16}: color_data = 12'haaa;
			{8'd108, 8'd17}: color_data = 12'h999;
			{8'd108, 8'd18}: color_data = 12'h999;
			{8'd108, 8'd19}: color_data = 12'h999;
			{8'd108, 8'd20}: color_data = 12'h999;
			{8'd108, 8'd21}: color_data = 12'h999;
			{8'd108, 8'd22}: color_data = 12'h999;
			{8'd108, 8'd23}: color_data = 12'h999;
			{8'd108, 8'd24}: color_data = 12'h999;
			{8'd108, 8'd25}: color_data = 12'h999;
			{8'd108, 8'd26}: color_data = 12'h999;
			{8'd108, 8'd27}: color_data = 12'h999;
			{8'd108, 8'd28}: color_data = 12'h999;
			{8'd108, 8'd29}: color_data = 12'h899;
			{8'd108, 8'd30}: color_data = 12'h7aa;
			{8'd108, 8'd31}: color_data = 12'hc11;
			{8'd108, 8'd32}: color_data = 12'hd21;
			{8'd108, 8'd33}: color_data = 12'hd31;
			{8'd108, 8'd34}: color_data = 12'hd31;
			{8'd108, 8'd35}: color_data = 12'hd41;
			{8'd108, 8'd36}: color_data = 12'he41;
			{8'd108, 8'd37}: color_data = 12'hd41;
			{8'd108, 8'd38}: color_data = 12'hd40;
			{8'd108, 8'd39}: color_data = 12'h799;
			{8'd108, 8'd40}: color_data = 12'h788;
			{8'd108, 8'd41}: color_data = 12'h788;
			{8'd108, 8'd42}: color_data = 12'h788;
			{8'd108, 8'd43}: color_data = 12'h788;
			{8'd108, 8'd44}: color_data = 12'h788;
			{8'd108, 8'd46}: color_data = 12'hd70;
			{8'd108, 8'd47}: color_data = 12'he80;
			{8'd108, 8'd48}: color_data = 12'he90;
			{8'd108, 8'd49}: color_data = 12'he90;
			{8'd108, 8'd50}: color_data = 12'he90;
			{8'd108, 8'd51}: color_data = 12'hd90;
			{8'd108, 8'd52}: color_data = 12'hc80;
			{8'd108, 8'd53}: color_data = 12'h677;
			{8'd108, 8'd54}: color_data = 12'h777;
			{8'd108, 8'd55}: color_data = 12'h777;
			{8'd108, 8'd56}: color_data = 12'h666;
			{8'd108, 8'd57}: color_data = 12'h666;
			{8'd108, 8'd58}: color_data = 12'h666;
			{8'd108, 8'd59}: color_data = 12'h666;
			{8'd108, 8'd60}: color_data = 12'h666;
			{8'd108, 8'd61}: color_data = 12'h666;
			{8'd108, 8'd62}: color_data = 12'h666;
			{8'd108, 8'd63}: color_data = 12'h666;
			{8'd108, 8'd64}: color_data = 12'h666;
			{8'd108, 8'd65}: color_data = 12'h666;
			{8'd108, 8'd66}: color_data = 12'h666;
			{8'd108, 8'd67}: color_data = 12'h666;
			{8'd108, 8'd68}: color_data = 12'h666;
			{8'd108, 8'd69}: color_data = 12'h555;
			{8'd108, 8'd70}: color_data = 12'h555;
			{8'd108, 8'd71}: color_data = 12'h555;
			{8'd108, 8'd72}: color_data = 12'h555;
			{8'd108, 8'd73}: color_data = 12'h555;
			{8'd108, 8'd74}: color_data = 12'h555;
			{8'd108, 8'd75}: color_data = 12'h555;
			{8'd108, 8'd76}: color_data = 12'h555;
			{8'd108, 8'd77}: color_data = 12'h555;
			{8'd108, 8'd78}: color_data = 12'h555;
			{8'd108, 8'd79}: color_data = 12'h555;
			{8'd108, 8'd80}: color_data = 12'h555;
			{8'd108, 8'd81}: color_data = 12'h555;
			{8'd108, 8'd82}: color_data = 12'h444;
			{8'd108, 8'd83}: color_data = 12'h444;
			{8'd108, 8'd84}: color_data = 12'h444;
			{8'd108, 8'd85}: color_data = 12'h444;
			{8'd108, 8'd86}: color_data = 12'h444;
			{8'd108, 8'd87}: color_data = 12'h444;
			{8'd108, 8'd88}: color_data = 12'h444;
			{8'd108, 8'd89}: color_data = 12'h444;
			{8'd108, 8'd90}: color_data = 12'h444;
			{8'd108, 8'd91}: color_data = 12'h444;
			{8'd108, 8'd92}: color_data = 12'h444;
			{8'd108, 8'd93}: color_data = 12'h444;
			{8'd108, 8'd94}: color_data = 12'h444;
			{8'd108, 8'd95}: color_data = 12'h333;
			{8'd108, 8'd96}: color_data = 12'h333;
			{8'd108, 8'd97}: color_data = 12'h333;
			{8'd108, 8'd98}: color_data = 12'h333;
			{8'd108, 8'd99}: color_data = 12'h333;
			{8'd108, 8'd100}: color_data = 12'h333;
			{8'd108, 8'd101}: color_data = 12'h333;
			{8'd108, 8'd102}: color_data = 12'h333;
			{8'd108, 8'd103}: color_data = 12'h333;
			{8'd108, 8'd104}: color_data = 12'h333;
			{8'd108, 8'd105}: color_data = 12'h333;
			{8'd108, 8'd106}: color_data = 12'h333;
			{8'd108, 8'd107}: color_data = 12'h333;
			{8'd108, 8'd108}: color_data = 12'h222;
			{8'd108, 8'd109}: color_data = 12'h222;
			{8'd108, 8'd110}: color_data = 12'h222;
			{8'd108, 8'd111}: color_data = 12'h222;
			{8'd108, 8'd112}: color_data = 12'h222;
			{8'd108, 8'd113}: color_data = 12'h222;
			{8'd108, 8'd114}: color_data = 12'h222;
			{8'd108, 8'd115}: color_data = 12'h222;
			{8'd108, 8'd116}: color_data = 12'h222;
			{8'd108, 8'd117}: color_data = 12'h222;
			{8'd108, 8'd118}: color_data = 12'h222;
			{8'd108, 8'd119}: color_data = 12'h222;
			{8'd108, 8'd120}: color_data = 12'h222;
			{8'd108, 8'd121}: color_data = 12'h111;
			{8'd108, 8'd122}: color_data = 12'h444;
			{8'd108, 8'd123}: color_data = 12'hddd;
			{8'd108, 8'd124}: color_data = 12'hfff;
			{8'd108, 8'd125}: color_data = 12'h777;
			{8'd108, 8'd126}: color_data = 12'h432;
			{8'd108, 8'd127}: color_data = 12'h642;
			{8'd108, 8'd128}: color_data = 12'h532;
			{8'd108, 8'd129}: color_data = 12'h632;
			{8'd108, 8'd130}: color_data = 12'h654;
			{8'd108, 8'd131}: color_data = 12'heee;
			{8'd108, 8'd132}: color_data = 12'hfff;
			{8'd108, 8'd133}: color_data = 12'hfff;
			{8'd108, 8'd134}: color_data = 12'hfff;
			{8'd108, 8'd135}: color_data = 12'hfff;
			{8'd108, 8'd136}: color_data = 12'hfff;
			{8'd108, 8'd137}: color_data = 12'hfff;
			{8'd108, 8'd138}: color_data = 12'hfff;
			{8'd108, 8'd139}: color_data = 12'hfff;
			{8'd108, 8'd140}: color_data = 12'hddd;
			{8'd108, 8'd141}: color_data = 12'hccc;
			{8'd109, 8'd0}: color_data = 12'hbbb;
			{8'd109, 8'd1}: color_data = 12'hbbb;
			{8'd109, 8'd2}: color_data = 12'hbbb;
			{8'd109, 8'd3}: color_data = 12'hbbb;
			{8'd109, 8'd4}: color_data = 12'haaa;
			{8'd109, 8'd5}: color_data = 12'haaa;
			{8'd109, 8'd6}: color_data = 12'haaa;
			{8'd109, 8'd7}: color_data = 12'haaa;
			{8'd109, 8'd8}: color_data = 12'haaa;
			{8'd109, 8'd9}: color_data = 12'haaa;
			{8'd109, 8'd10}: color_data = 12'haaa;
			{8'd109, 8'd11}: color_data = 12'haaa;
			{8'd109, 8'd12}: color_data = 12'haaa;
			{8'd109, 8'd13}: color_data = 12'haaa;
			{8'd109, 8'd14}: color_data = 12'haaa;
			{8'd109, 8'd15}: color_data = 12'haaa;
			{8'd109, 8'd16}: color_data = 12'haaa;
			{8'd109, 8'd17}: color_data = 12'h999;
			{8'd109, 8'd18}: color_data = 12'h999;
			{8'd109, 8'd19}: color_data = 12'h999;
			{8'd109, 8'd20}: color_data = 12'h999;
			{8'd109, 8'd21}: color_data = 12'h999;
			{8'd109, 8'd22}: color_data = 12'h999;
			{8'd109, 8'd23}: color_data = 12'h999;
			{8'd109, 8'd24}: color_data = 12'h999;
			{8'd109, 8'd25}: color_data = 12'h999;
			{8'd109, 8'd26}: color_data = 12'h999;
			{8'd109, 8'd27}: color_data = 12'h999;
			{8'd109, 8'd28}: color_data = 12'h999;
			{8'd109, 8'd29}: color_data = 12'h999;
			{8'd109, 8'd30}: color_data = 12'hc00;
			{8'd109, 8'd31}: color_data = 12'hd21;
			{8'd109, 8'd32}: color_data = 12'he21;
			{8'd109, 8'd33}: color_data = 12'hd31;
			{8'd109, 8'd34}: color_data = 12'hd31;
			{8'd109, 8'd35}: color_data = 12'he41;
			{8'd109, 8'd36}: color_data = 12'he41;
			{8'd109, 8'd37}: color_data = 12'hd41;
			{8'd109, 8'd38}: color_data = 12'he40;
			{8'd109, 8'd39}: color_data = 12'h788;
			{8'd109, 8'd40}: color_data = 12'h888;
			{8'd109, 8'd41}: color_data = 12'h888;
			{8'd109, 8'd42}: color_data = 12'h888;
			{8'd109, 8'd43}: color_data = 12'h888;
			{8'd109, 8'd44}: color_data = 12'h777;
			{8'd109, 8'd45}: color_data = 12'h679;
			{8'd109, 8'd46}: color_data = 12'hd70;
			{8'd109, 8'd47}: color_data = 12'hd80;
			{8'd109, 8'd48}: color_data = 12'hd80;
			{8'd109, 8'd49}: color_data = 12'hd80;
			{8'd109, 8'd50}: color_data = 12'hd90;
			{8'd109, 8'd51}: color_data = 12'hc80;
			{8'd109, 8'd52}: color_data = 12'hb70;
			{8'd109, 8'd53}: color_data = 12'h667;
			{8'd109, 8'd54}: color_data = 12'h777;
			{8'd109, 8'd55}: color_data = 12'h777;
			{8'd109, 8'd56}: color_data = 12'h666;
			{8'd109, 8'd57}: color_data = 12'h666;
			{8'd109, 8'd58}: color_data = 12'h666;
			{8'd109, 8'd59}: color_data = 12'h666;
			{8'd109, 8'd60}: color_data = 12'h666;
			{8'd109, 8'd61}: color_data = 12'h666;
			{8'd109, 8'd62}: color_data = 12'h666;
			{8'd109, 8'd63}: color_data = 12'h666;
			{8'd109, 8'd64}: color_data = 12'h666;
			{8'd109, 8'd65}: color_data = 12'h666;
			{8'd109, 8'd66}: color_data = 12'h666;
			{8'd109, 8'd67}: color_data = 12'h666;
			{8'd109, 8'd68}: color_data = 12'h666;
			{8'd109, 8'd69}: color_data = 12'h555;
			{8'd109, 8'd70}: color_data = 12'h555;
			{8'd109, 8'd71}: color_data = 12'h555;
			{8'd109, 8'd72}: color_data = 12'h555;
			{8'd109, 8'd73}: color_data = 12'h555;
			{8'd109, 8'd74}: color_data = 12'h555;
			{8'd109, 8'd75}: color_data = 12'h555;
			{8'd109, 8'd76}: color_data = 12'h555;
			{8'd109, 8'd77}: color_data = 12'h555;
			{8'd109, 8'd78}: color_data = 12'h555;
			{8'd109, 8'd79}: color_data = 12'h555;
			{8'd109, 8'd80}: color_data = 12'h555;
			{8'd109, 8'd81}: color_data = 12'h555;
			{8'd109, 8'd82}: color_data = 12'h444;
			{8'd109, 8'd83}: color_data = 12'h444;
			{8'd109, 8'd84}: color_data = 12'h444;
			{8'd109, 8'd85}: color_data = 12'h444;
			{8'd109, 8'd86}: color_data = 12'h444;
			{8'd109, 8'd87}: color_data = 12'h444;
			{8'd109, 8'd88}: color_data = 12'h444;
			{8'd109, 8'd89}: color_data = 12'h444;
			{8'd109, 8'd90}: color_data = 12'h444;
			{8'd109, 8'd91}: color_data = 12'h444;
			{8'd109, 8'd92}: color_data = 12'h444;
			{8'd109, 8'd93}: color_data = 12'h444;
			{8'd109, 8'd94}: color_data = 12'h444;
			{8'd109, 8'd95}: color_data = 12'h333;
			{8'd109, 8'd96}: color_data = 12'h333;
			{8'd109, 8'd97}: color_data = 12'h333;
			{8'd109, 8'd98}: color_data = 12'h333;
			{8'd109, 8'd99}: color_data = 12'h333;
			{8'd109, 8'd100}: color_data = 12'h333;
			{8'd109, 8'd101}: color_data = 12'h333;
			{8'd109, 8'd102}: color_data = 12'h333;
			{8'd109, 8'd103}: color_data = 12'h333;
			{8'd109, 8'd104}: color_data = 12'h333;
			{8'd109, 8'd105}: color_data = 12'h333;
			{8'd109, 8'd106}: color_data = 12'h333;
			{8'd109, 8'd107}: color_data = 12'h333;
			{8'd109, 8'd108}: color_data = 12'h222;
			{8'd109, 8'd109}: color_data = 12'h222;
			{8'd109, 8'd110}: color_data = 12'h222;
			{8'd109, 8'd111}: color_data = 12'h222;
			{8'd109, 8'd112}: color_data = 12'h222;
			{8'd109, 8'd113}: color_data = 12'h222;
			{8'd109, 8'd114}: color_data = 12'h222;
			{8'd109, 8'd115}: color_data = 12'h222;
			{8'd109, 8'd116}: color_data = 12'h222;
			{8'd109, 8'd117}: color_data = 12'h222;
			{8'd109, 8'd118}: color_data = 12'h222;
			{8'd109, 8'd119}: color_data = 12'h222;
			{8'd109, 8'd120}: color_data = 12'h222;
			{8'd109, 8'd121}: color_data = 12'h111;
			{8'd109, 8'd122}: color_data = 12'h444;
			{8'd109, 8'd123}: color_data = 12'hddd;
			{8'd109, 8'd124}: color_data = 12'hddd;
			{8'd109, 8'd125}: color_data = 12'h433;
			{8'd109, 8'd126}: color_data = 12'h642;
			{8'd109, 8'd127}: color_data = 12'h432;
			{8'd109, 8'd128}: color_data = 12'h532;
			{8'd109, 8'd129}: color_data = 12'h852;
			{8'd109, 8'd130}: color_data = 12'h654;
			{8'd109, 8'd131}: color_data = 12'hdee;
			{8'd109, 8'd132}: color_data = 12'hfff;
			{8'd109, 8'd133}: color_data = 12'hfff;
			{8'd109, 8'd134}: color_data = 12'hfff;
			{8'd109, 8'd135}: color_data = 12'hfff;
			{8'd109, 8'd136}: color_data = 12'hfff;
			{8'd109, 8'd137}: color_data = 12'hfff;
			{8'd109, 8'd138}: color_data = 12'hfff;
			{8'd109, 8'd139}: color_data = 12'hfff;
			{8'd109, 8'd140}: color_data = 12'hddd;
			{8'd109, 8'd141}: color_data = 12'hddd;
			{8'd110, 8'd0}: color_data = 12'hbbb;
			{8'd110, 8'd1}: color_data = 12'hbbb;
			{8'd110, 8'd2}: color_data = 12'hbbb;
			{8'd110, 8'd3}: color_data = 12'hbbb;
			{8'd110, 8'd4}: color_data = 12'haaa;
			{8'd110, 8'd5}: color_data = 12'haaa;
			{8'd110, 8'd6}: color_data = 12'haaa;
			{8'd110, 8'd7}: color_data = 12'haaa;
			{8'd110, 8'd8}: color_data = 12'haaa;
			{8'd110, 8'd9}: color_data = 12'haaa;
			{8'd110, 8'd10}: color_data = 12'haaa;
			{8'd110, 8'd11}: color_data = 12'haaa;
			{8'd110, 8'd12}: color_data = 12'haaa;
			{8'd110, 8'd13}: color_data = 12'haaa;
			{8'd110, 8'd14}: color_data = 12'haaa;
			{8'd110, 8'd15}: color_data = 12'haaa;
			{8'd110, 8'd16}: color_data = 12'h999;
			{8'd110, 8'd17}: color_data = 12'h999;
			{8'd110, 8'd18}: color_data = 12'h999;
			{8'd110, 8'd19}: color_data = 12'h999;
			{8'd110, 8'd20}: color_data = 12'h999;
			{8'd110, 8'd21}: color_data = 12'h999;
			{8'd110, 8'd22}: color_data = 12'h999;
			{8'd110, 8'd23}: color_data = 12'h999;
			{8'd110, 8'd24}: color_data = 12'h999;
			{8'd110, 8'd25}: color_data = 12'h999;
			{8'd110, 8'd26}: color_data = 12'h999;
			{8'd110, 8'd27}: color_data = 12'h999;
			{8'd110, 8'd28}: color_data = 12'h999;
			{8'd110, 8'd29}: color_data = 12'h899;
			{8'd110, 8'd30}: color_data = 12'hf00;
			{8'd110, 8'd31}: color_data = 12'hd21;
			{8'd110, 8'd32}: color_data = 12'he21;
			{8'd110, 8'd33}: color_data = 12'hd31;
			{8'd110, 8'd34}: color_data = 12'he31;
			{8'd110, 8'd35}: color_data = 12'he41;
			{8'd110, 8'd36}: color_data = 12'he41;
			{8'd110, 8'd37}: color_data = 12'hd41;
			{8'd110, 8'd38}: color_data = 12'he30;
			{8'd110, 8'd39}: color_data = 12'h788;
			{8'd110, 8'd40}: color_data = 12'h888;
			{8'd110, 8'd41}: color_data = 12'h888;
			{8'd110, 8'd42}: color_data = 12'h888;
			{8'd110, 8'd43}: color_data = 12'h888;
			{8'd110, 8'd44}: color_data = 12'h888;
			{8'd110, 8'd45}: color_data = 12'h777;
			{8'd110, 8'd47}: color_data = 12'hb60;
			{8'd110, 8'd48}: color_data = 12'hb70;
			{8'd110, 8'd49}: color_data = 12'hb70;
			{8'd110, 8'd50}: color_data = 12'hb70;
			{8'd110, 8'd51}: color_data = 12'hb70;
			{8'd110, 8'd53}: color_data = 12'h667;
			{8'd110, 8'd54}: color_data = 12'h777;
			{8'd110, 8'd55}: color_data = 12'h777;
			{8'd110, 8'd56}: color_data = 12'h666;
			{8'd110, 8'd57}: color_data = 12'h666;
			{8'd110, 8'd58}: color_data = 12'h666;
			{8'd110, 8'd59}: color_data = 12'h666;
			{8'd110, 8'd60}: color_data = 12'h666;
			{8'd110, 8'd61}: color_data = 12'h666;
			{8'd110, 8'd62}: color_data = 12'h666;
			{8'd110, 8'd63}: color_data = 12'h666;
			{8'd110, 8'd64}: color_data = 12'h666;
			{8'd110, 8'd65}: color_data = 12'h666;
			{8'd110, 8'd66}: color_data = 12'h666;
			{8'd110, 8'd67}: color_data = 12'h666;
			{8'd110, 8'd68}: color_data = 12'h666;
			{8'd110, 8'd69}: color_data = 12'h555;
			{8'd110, 8'd70}: color_data = 12'h555;
			{8'd110, 8'd71}: color_data = 12'h555;
			{8'd110, 8'd72}: color_data = 12'h555;
			{8'd110, 8'd73}: color_data = 12'h555;
			{8'd110, 8'd74}: color_data = 12'h555;
			{8'd110, 8'd75}: color_data = 12'h555;
			{8'd110, 8'd76}: color_data = 12'h555;
			{8'd110, 8'd77}: color_data = 12'h555;
			{8'd110, 8'd78}: color_data = 12'h555;
			{8'd110, 8'd79}: color_data = 12'h555;
			{8'd110, 8'd80}: color_data = 12'h555;
			{8'd110, 8'd81}: color_data = 12'h555;
			{8'd110, 8'd82}: color_data = 12'h444;
			{8'd110, 8'd83}: color_data = 12'h444;
			{8'd110, 8'd84}: color_data = 12'h444;
			{8'd110, 8'd85}: color_data = 12'h444;
			{8'd110, 8'd86}: color_data = 12'h444;
			{8'd110, 8'd87}: color_data = 12'h444;
			{8'd110, 8'd88}: color_data = 12'h444;
			{8'd110, 8'd89}: color_data = 12'h444;
			{8'd110, 8'd90}: color_data = 12'h444;
			{8'd110, 8'd91}: color_data = 12'h444;
			{8'd110, 8'd92}: color_data = 12'h444;
			{8'd110, 8'd93}: color_data = 12'h444;
			{8'd110, 8'd94}: color_data = 12'h444;
			{8'd110, 8'd95}: color_data = 12'h333;
			{8'd110, 8'd96}: color_data = 12'h333;
			{8'd110, 8'd97}: color_data = 12'h333;
			{8'd110, 8'd98}: color_data = 12'h333;
			{8'd110, 8'd99}: color_data = 12'h333;
			{8'd110, 8'd100}: color_data = 12'h333;
			{8'd110, 8'd101}: color_data = 12'h333;
			{8'd110, 8'd102}: color_data = 12'h333;
			{8'd110, 8'd103}: color_data = 12'h333;
			{8'd110, 8'd104}: color_data = 12'h333;
			{8'd110, 8'd105}: color_data = 12'h333;
			{8'd110, 8'd106}: color_data = 12'h333;
			{8'd110, 8'd107}: color_data = 12'h333;
			{8'd110, 8'd108}: color_data = 12'h222;
			{8'd110, 8'd109}: color_data = 12'h222;
			{8'd110, 8'd110}: color_data = 12'h222;
			{8'd110, 8'd111}: color_data = 12'h222;
			{8'd110, 8'd112}: color_data = 12'h222;
			{8'd110, 8'd113}: color_data = 12'h222;
			{8'd110, 8'd114}: color_data = 12'h222;
			{8'd110, 8'd115}: color_data = 12'h222;
			{8'd110, 8'd116}: color_data = 12'h222;
			{8'd110, 8'd117}: color_data = 12'h222;
			{8'd110, 8'd118}: color_data = 12'h222;
			{8'd110, 8'd119}: color_data = 12'h222;
			{8'd110, 8'd120}: color_data = 12'h222;
			{8'd110, 8'd121}: color_data = 12'h111;
			{8'd110, 8'd122}: color_data = 12'h555;
			{8'd110, 8'd123}: color_data = 12'heee;
			{8'd110, 8'd124}: color_data = 12'hdcc;
			{8'd110, 8'd125}: color_data = 12'h322;
			{8'd110, 8'd126}: color_data = 12'h532;
			{8'd110, 8'd127}: color_data = 12'h532;
			{8'd110, 8'd128}: color_data = 12'h432;
			{8'd110, 8'd129}: color_data = 12'h322;
			{8'd110, 8'd130}: color_data = 12'h444;
			{8'd110, 8'd131}: color_data = 12'hddd;
			{8'd110, 8'd132}: color_data = 12'hfff;
			{8'd110, 8'd133}: color_data = 12'hfff;
			{8'd110, 8'd134}: color_data = 12'hfff;
			{8'd110, 8'd135}: color_data = 12'hfff;
			{8'd110, 8'd136}: color_data = 12'hfff;
			{8'd110, 8'd137}: color_data = 12'hfff;
			{8'd110, 8'd138}: color_data = 12'hfff;
			{8'd110, 8'd139}: color_data = 12'hfff;
			{8'd110, 8'd140}: color_data = 12'heee;
			{8'd110, 8'd141}: color_data = 12'hddd;
			{8'd111, 8'd0}: color_data = 12'hbbb;
			{8'd111, 8'd1}: color_data = 12'hbbb;
			{8'd111, 8'd2}: color_data = 12'hbbb;
			{8'd111, 8'd3}: color_data = 12'hbbb;
			{8'd111, 8'd4}: color_data = 12'haaa;
			{8'd111, 8'd5}: color_data = 12'haaa;
			{8'd111, 8'd6}: color_data = 12'haaa;
			{8'd111, 8'd7}: color_data = 12'haaa;
			{8'd111, 8'd8}: color_data = 12'haaa;
			{8'd111, 8'd9}: color_data = 12'haaa;
			{8'd111, 8'd10}: color_data = 12'haaa;
			{8'd111, 8'd11}: color_data = 12'haaa;
			{8'd111, 8'd12}: color_data = 12'haaa;
			{8'd111, 8'd13}: color_data = 12'haaa;
			{8'd111, 8'd14}: color_data = 12'haaa;
			{8'd111, 8'd15}: color_data = 12'haaa;
			{8'd111, 8'd16}: color_data = 12'h999;
			{8'd111, 8'd17}: color_data = 12'h999;
			{8'd111, 8'd18}: color_data = 12'h999;
			{8'd111, 8'd19}: color_data = 12'h999;
			{8'd111, 8'd20}: color_data = 12'h999;
			{8'd111, 8'd21}: color_data = 12'h999;
			{8'd111, 8'd22}: color_data = 12'h999;
			{8'd111, 8'd23}: color_data = 12'h999;
			{8'd111, 8'd24}: color_data = 12'h999;
			{8'd111, 8'd25}: color_data = 12'h999;
			{8'd111, 8'd26}: color_data = 12'h999;
			{8'd111, 8'd27}: color_data = 12'h999;
			{8'd111, 8'd28}: color_data = 12'h999;
			{8'd111, 8'd29}: color_data = 12'h888;
			{8'd111, 8'd31}: color_data = 12'hd11;
			{8'd111, 8'd32}: color_data = 12'hd21;
			{8'd111, 8'd33}: color_data = 12'hd21;
			{8'd111, 8'd34}: color_data = 12'hd31;
			{8'd111, 8'd35}: color_data = 12'hd31;
			{8'd111, 8'd36}: color_data = 12'hd41;
			{8'd111, 8'd37}: color_data = 12'hd41;
			{8'd111, 8'd39}: color_data = 12'h888;
			{8'd111, 8'd40}: color_data = 12'h888;
			{8'd111, 8'd41}: color_data = 12'h888;
			{8'd111, 8'd42}: color_data = 12'h888;
			{8'd111, 8'd43}: color_data = 12'h777;
			{8'd111, 8'd44}: color_data = 12'h777;
			{8'd111, 8'd45}: color_data = 12'h777;
			{8'd111, 8'd46}: color_data = 12'h777;
			{8'd111, 8'd47}: color_data = 12'h778;
			{8'd111, 8'd48}: color_data = 12'h677;
			{8'd111, 8'd49}: color_data = 12'h777;
			{8'd111, 8'd50}: color_data = 12'h677;
			{8'd111, 8'd51}: color_data = 12'h45a;
			{8'd111, 8'd52}: color_data = 12'h666;
			{8'd111, 8'd53}: color_data = 12'h666;
			{8'd111, 8'd54}: color_data = 12'h777;
			{8'd111, 8'd55}: color_data = 12'h777;
			{8'd111, 8'd56}: color_data = 12'h666;
			{8'd111, 8'd57}: color_data = 12'h666;
			{8'd111, 8'd58}: color_data = 12'h666;
			{8'd111, 8'd59}: color_data = 12'h666;
			{8'd111, 8'd60}: color_data = 12'h666;
			{8'd111, 8'd61}: color_data = 12'h666;
			{8'd111, 8'd62}: color_data = 12'h666;
			{8'd111, 8'd63}: color_data = 12'h666;
			{8'd111, 8'd64}: color_data = 12'h666;
			{8'd111, 8'd65}: color_data = 12'h666;
			{8'd111, 8'd66}: color_data = 12'h666;
			{8'd111, 8'd67}: color_data = 12'h666;
			{8'd111, 8'd68}: color_data = 12'h666;
			{8'd111, 8'd69}: color_data = 12'h555;
			{8'd111, 8'd70}: color_data = 12'h555;
			{8'd111, 8'd71}: color_data = 12'h555;
			{8'd111, 8'd72}: color_data = 12'h555;
			{8'd111, 8'd73}: color_data = 12'h555;
			{8'd111, 8'd74}: color_data = 12'h555;
			{8'd111, 8'd75}: color_data = 12'h555;
			{8'd111, 8'd76}: color_data = 12'h555;
			{8'd111, 8'd77}: color_data = 12'h555;
			{8'd111, 8'd78}: color_data = 12'h555;
			{8'd111, 8'd79}: color_data = 12'h555;
			{8'd111, 8'd80}: color_data = 12'h555;
			{8'd111, 8'd81}: color_data = 12'h555;
			{8'd111, 8'd82}: color_data = 12'h444;
			{8'd111, 8'd83}: color_data = 12'h444;
			{8'd111, 8'd84}: color_data = 12'h444;
			{8'd111, 8'd85}: color_data = 12'h444;
			{8'd111, 8'd86}: color_data = 12'h444;
			{8'd111, 8'd87}: color_data = 12'h444;
			{8'd111, 8'd88}: color_data = 12'h444;
			{8'd111, 8'd89}: color_data = 12'h444;
			{8'd111, 8'd90}: color_data = 12'h444;
			{8'd111, 8'd91}: color_data = 12'h444;
			{8'd111, 8'd92}: color_data = 12'h444;
			{8'd111, 8'd93}: color_data = 12'h444;
			{8'd111, 8'd94}: color_data = 12'h444;
			{8'd111, 8'd95}: color_data = 12'h333;
			{8'd111, 8'd96}: color_data = 12'h333;
			{8'd111, 8'd97}: color_data = 12'h333;
			{8'd111, 8'd98}: color_data = 12'h333;
			{8'd111, 8'd99}: color_data = 12'h333;
			{8'd111, 8'd100}: color_data = 12'h333;
			{8'd111, 8'd101}: color_data = 12'h333;
			{8'd111, 8'd102}: color_data = 12'h333;
			{8'd111, 8'd103}: color_data = 12'h333;
			{8'd111, 8'd104}: color_data = 12'h333;
			{8'd111, 8'd105}: color_data = 12'h333;
			{8'd111, 8'd106}: color_data = 12'h333;
			{8'd111, 8'd107}: color_data = 12'h333;
			{8'd111, 8'd108}: color_data = 12'h222;
			{8'd111, 8'd109}: color_data = 12'h222;
			{8'd111, 8'd110}: color_data = 12'h222;
			{8'd111, 8'd111}: color_data = 12'h222;
			{8'd111, 8'd112}: color_data = 12'h222;
			{8'd111, 8'd113}: color_data = 12'h222;
			{8'd111, 8'd114}: color_data = 12'h222;
			{8'd111, 8'd115}: color_data = 12'h222;
			{8'd111, 8'd116}: color_data = 12'h222;
			{8'd111, 8'd117}: color_data = 12'h222;
			{8'd111, 8'd118}: color_data = 12'h222;
			{8'd111, 8'd119}: color_data = 12'h222;
			{8'd111, 8'd120}: color_data = 12'h222;
			{8'd111, 8'd121}: color_data = 12'h111;
			{8'd111, 8'd122}: color_data = 12'h666;
			{8'd111, 8'd123}: color_data = 12'hddd;
			{8'd111, 8'd124}: color_data = 12'h877;
			{8'd111, 8'd125}: color_data = 12'h334;
			{8'd111, 8'd126}: color_data = 12'h338;
			{8'd111, 8'd127}: color_data = 12'h338;
			{8'd111, 8'd128}: color_data = 12'h338;
			{8'd111, 8'd129}: color_data = 12'h225;
			{8'd111, 8'd130}: color_data = 12'h444;
			{8'd111, 8'd131}: color_data = 12'hccc;
			{8'd111, 8'd132}: color_data = 12'heee;
			{8'd111, 8'd133}: color_data = 12'hfff;
			{8'd111, 8'd134}: color_data = 12'hfff;
			{8'd111, 8'd135}: color_data = 12'hfff;
			{8'd111, 8'd136}: color_data = 12'hfff;
			{8'd111, 8'd137}: color_data = 12'hfff;
			{8'd111, 8'd138}: color_data = 12'hfff;
			{8'd111, 8'd139}: color_data = 12'hfff;
			{8'd111, 8'd140}: color_data = 12'heee;
			{8'd111, 8'd141}: color_data = 12'hddd;
			{8'd112, 8'd0}: color_data = 12'hbbb;
			{8'd112, 8'd1}: color_data = 12'hbbb;
			{8'd112, 8'd2}: color_data = 12'hbbb;
			{8'd112, 8'd3}: color_data = 12'hbbb;
			{8'd112, 8'd4}: color_data = 12'haaa;
			{8'd112, 8'd5}: color_data = 12'haaa;
			{8'd112, 8'd6}: color_data = 12'haaa;
			{8'd112, 8'd7}: color_data = 12'haaa;
			{8'd112, 8'd8}: color_data = 12'haaa;
			{8'd112, 8'd9}: color_data = 12'haaa;
			{8'd112, 8'd10}: color_data = 12'haaa;
			{8'd112, 8'd11}: color_data = 12'haaa;
			{8'd112, 8'd12}: color_data = 12'haaa;
			{8'd112, 8'd13}: color_data = 12'haaa;
			{8'd112, 8'd14}: color_data = 12'haaa;
			{8'd112, 8'd15}: color_data = 12'haaa;
			{8'd112, 8'd16}: color_data = 12'h999;
			{8'd112, 8'd17}: color_data = 12'h999;
			{8'd112, 8'd18}: color_data = 12'h999;
			{8'd112, 8'd19}: color_data = 12'h999;
			{8'd112, 8'd20}: color_data = 12'h999;
			{8'd112, 8'd21}: color_data = 12'h999;
			{8'd112, 8'd22}: color_data = 12'h999;
			{8'd112, 8'd23}: color_data = 12'h999;
			{8'd112, 8'd24}: color_data = 12'h999;
			{8'd112, 8'd25}: color_data = 12'h999;
			{8'd112, 8'd26}: color_data = 12'h999;
			{8'd112, 8'd27}: color_data = 12'h999;
			{8'd112, 8'd28}: color_data = 12'h999;
			{8'd112, 8'd29}: color_data = 12'h888;
			{8'd112, 8'd30}: color_data = 12'h0ff;
			{8'd112, 8'd31}: color_data = 12'h7aa;
			{8'd112, 8'd32}: color_data = 12'ha66;
			{8'd112, 8'd33}: color_data = 12'h976;
			{8'd112, 8'd34}: color_data = 12'h69b;
			{8'd112, 8'd35}: color_data = 12'h777;
			{8'd112, 8'd36}: color_data = 12'ha65;
			{8'd112, 8'd37}: color_data = 12'h778;
			{8'd112, 8'd38}: color_data = 12'h777;
			{8'd112, 8'd39}: color_data = 12'h888;
			{8'd112, 8'd40}: color_data = 12'h888;
			{8'd112, 8'd41}: color_data = 12'h888;
			{8'd112, 8'd42}: color_data = 12'h888;
			{8'd112, 8'd43}: color_data = 12'h777;
			{8'd112, 8'd44}: color_data = 12'h777;
			{8'd112, 8'd45}: color_data = 12'h777;
			{8'd112, 8'd46}: color_data = 12'h777;
			{8'd112, 8'd47}: color_data = 12'h777;
			{8'd112, 8'd48}: color_data = 12'h777;
			{8'd112, 8'd49}: color_data = 12'h777;
			{8'd112, 8'd50}: color_data = 12'h777;
			{8'd112, 8'd51}: color_data = 12'h777;
			{8'd112, 8'd52}: color_data = 12'h777;
			{8'd112, 8'd53}: color_data = 12'h777;
			{8'd112, 8'd54}: color_data = 12'h777;
			{8'd112, 8'd55}: color_data = 12'h777;
			{8'd112, 8'd56}: color_data = 12'h666;
			{8'd112, 8'd57}: color_data = 12'h666;
			{8'd112, 8'd58}: color_data = 12'h666;
			{8'd112, 8'd59}: color_data = 12'h666;
			{8'd112, 8'd60}: color_data = 12'h666;
			{8'd112, 8'd61}: color_data = 12'h666;
			{8'd112, 8'd62}: color_data = 12'h666;
			{8'd112, 8'd63}: color_data = 12'h666;
			{8'd112, 8'd64}: color_data = 12'h666;
			{8'd112, 8'd65}: color_data = 12'h666;
			{8'd112, 8'd66}: color_data = 12'h666;
			{8'd112, 8'd67}: color_data = 12'h666;
			{8'd112, 8'd68}: color_data = 12'h666;
			{8'd112, 8'd69}: color_data = 12'h555;
			{8'd112, 8'd70}: color_data = 12'h555;
			{8'd112, 8'd71}: color_data = 12'h555;
			{8'd112, 8'd72}: color_data = 12'h555;
			{8'd112, 8'd73}: color_data = 12'h555;
			{8'd112, 8'd74}: color_data = 12'h555;
			{8'd112, 8'd75}: color_data = 12'h555;
			{8'd112, 8'd76}: color_data = 12'h555;
			{8'd112, 8'd77}: color_data = 12'h555;
			{8'd112, 8'd78}: color_data = 12'h555;
			{8'd112, 8'd79}: color_data = 12'h555;
			{8'd112, 8'd80}: color_data = 12'h555;
			{8'd112, 8'd81}: color_data = 12'h555;
			{8'd112, 8'd82}: color_data = 12'h444;
			{8'd112, 8'd83}: color_data = 12'h444;
			{8'd112, 8'd84}: color_data = 12'h444;
			{8'd112, 8'd85}: color_data = 12'h444;
			{8'd112, 8'd86}: color_data = 12'h444;
			{8'd112, 8'd87}: color_data = 12'h444;
			{8'd112, 8'd88}: color_data = 12'h444;
			{8'd112, 8'd89}: color_data = 12'h444;
			{8'd112, 8'd90}: color_data = 12'h444;
			{8'd112, 8'd91}: color_data = 12'h444;
			{8'd112, 8'd92}: color_data = 12'h444;
			{8'd112, 8'd93}: color_data = 12'h444;
			{8'd112, 8'd94}: color_data = 12'h444;
			{8'd112, 8'd95}: color_data = 12'h333;
			{8'd112, 8'd96}: color_data = 12'h333;
			{8'd112, 8'd97}: color_data = 12'h333;
			{8'd112, 8'd98}: color_data = 12'h333;
			{8'd112, 8'd99}: color_data = 12'h333;
			{8'd112, 8'd100}: color_data = 12'h333;
			{8'd112, 8'd101}: color_data = 12'h333;
			{8'd112, 8'd102}: color_data = 12'h333;
			{8'd112, 8'd103}: color_data = 12'h333;
			{8'd112, 8'd104}: color_data = 12'h333;
			{8'd112, 8'd105}: color_data = 12'h333;
			{8'd112, 8'd106}: color_data = 12'h333;
			{8'd112, 8'd107}: color_data = 12'h333;
			{8'd112, 8'd108}: color_data = 12'h222;
			{8'd112, 8'd109}: color_data = 12'h222;
			{8'd112, 8'd110}: color_data = 12'h222;
			{8'd112, 8'd111}: color_data = 12'h222;
			{8'd112, 8'd112}: color_data = 12'h222;
			{8'd112, 8'd113}: color_data = 12'h222;
			{8'd112, 8'd114}: color_data = 12'h222;
			{8'd112, 8'd115}: color_data = 12'h222;
			{8'd112, 8'd116}: color_data = 12'h222;
			{8'd112, 8'd117}: color_data = 12'h222;
			{8'd112, 8'd118}: color_data = 12'h222;
			{8'd112, 8'd119}: color_data = 12'h222;
			{8'd112, 8'd120}: color_data = 12'h222;
			{8'd112, 8'd121}: color_data = 12'h222;
			{8'd112, 8'd122}: color_data = 12'h666;
			{8'd112, 8'd123}: color_data = 12'h766;
			{8'd112, 8'd124}: color_data = 12'h336;
			{8'd112, 8'd125}: color_data = 12'h34c;
			{8'd112, 8'd126}: color_data = 12'h34d;
			{8'd112, 8'd127}: color_data = 12'h44b;
			{8'd112, 8'd128}: color_data = 12'h569;
			{8'd112, 8'd129}: color_data = 12'h557;
			{8'd112, 8'd130}: color_data = 12'h555;
			{8'd112, 8'd131}: color_data = 12'hbbb;
			{8'd112, 8'd132}: color_data = 12'hddd;
			{8'd112, 8'd133}: color_data = 12'hfff;
			{8'd112, 8'd134}: color_data = 12'hfff;
			{8'd112, 8'd135}: color_data = 12'hfff;
			{8'd112, 8'd136}: color_data = 12'hfff;
			{8'd112, 8'd137}: color_data = 12'hfff;
			{8'd112, 8'd138}: color_data = 12'hfff;
			{8'd112, 8'd139}: color_data = 12'hfff;
			{8'd112, 8'd140}: color_data = 12'heee;
			{8'd112, 8'd141}: color_data = 12'heee;
			{8'd113, 8'd0}: color_data = 12'hbbb;
			{8'd113, 8'd1}: color_data = 12'hbbb;
			{8'd113, 8'd2}: color_data = 12'hbbb;
			{8'd113, 8'd3}: color_data = 12'hbbb;
			{8'd113, 8'd4}: color_data = 12'haaa;
			{8'd113, 8'd5}: color_data = 12'haaa;
			{8'd113, 8'd6}: color_data = 12'haaa;
			{8'd113, 8'd7}: color_data = 12'haaa;
			{8'd113, 8'd8}: color_data = 12'haaa;
			{8'd113, 8'd9}: color_data = 12'haaa;
			{8'd113, 8'd10}: color_data = 12'haaa;
			{8'd113, 8'd11}: color_data = 12'haaa;
			{8'd113, 8'd12}: color_data = 12'haaa;
			{8'd113, 8'd13}: color_data = 12'haaa;
			{8'd113, 8'd14}: color_data = 12'haaa;
			{8'd113, 8'd15}: color_data = 12'haaa;
			{8'd113, 8'd16}: color_data = 12'h999;
			{8'd113, 8'd17}: color_data = 12'h999;
			{8'd113, 8'd18}: color_data = 12'h999;
			{8'd113, 8'd19}: color_data = 12'h999;
			{8'd113, 8'd20}: color_data = 12'h999;
			{8'd113, 8'd21}: color_data = 12'h999;
			{8'd113, 8'd22}: color_data = 12'h999;
			{8'd113, 8'd23}: color_data = 12'h999;
			{8'd113, 8'd24}: color_data = 12'h999;
			{8'd113, 8'd25}: color_data = 12'h999;
			{8'd113, 8'd26}: color_data = 12'h999;
			{8'd113, 8'd27}: color_data = 12'h999;
			{8'd113, 8'd28}: color_data = 12'h888;
			{8'd113, 8'd29}: color_data = 12'h888;
			{8'd113, 8'd30}: color_data = 12'h888;
			{8'd113, 8'd31}: color_data = 12'h889;
			{8'd113, 8'd32}: color_data = 12'h888;
			{8'd113, 8'd33}: color_data = 12'h888;
			{8'd113, 8'd34}: color_data = 12'h888;
			{8'd113, 8'd35}: color_data = 12'h888;
			{8'd113, 8'd36}: color_data = 12'h888;
			{8'd113, 8'd37}: color_data = 12'h888;
			{8'd113, 8'd38}: color_data = 12'h888;
			{8'd113, 8'd39}: color_data = 12'h888;
			{8'd113, 8'd40}: color_data = 12'h888;
			{8'd113, 8'd41}: color_data = 12'h888;
			{8'd113, 8'd42}: color_data = 12'h888;
			{8'd113, 8'd43}: color_data = 12'h777;
			{8'd113, 8'd44}: color_data = 12'h777;
			{8'd113, 8'd45}: color_data = 12'h777;
			{8'd113, 8'd46}: color_data = 12'h777;
			{8'd113, 8'd47}: color_data = 12'h777;
			{8'd113, 8'd48}: color_data = 12'h777;
			{8'd113, 8'd49}: color_data = 12'h777;
			{8'd113, 8'd50}: color_data = 12'h777;
			{8'd113, 8'd51}: color_data = 12'h777;
			{8'd113, 8'd52}: color_data = 12'h777;
			{8'd113, 8'd53}: color_data = 12'h777;
			{8'd113, 8'd54}: color_data = 12'h777;
			{8'd113, 8'd55}: color_data = 12'h777;
			{8'd113, 8'd56}: color_data = 12'h666;
			{8'd113, 8'd57}: color_data = 12'h666;
			{8'd113, 8'd58}: color_data = 12'h666;
			{8'd113, 8'd59}: color_data = 12'h666;
			{8'd113, 8'd60}: color_data = 12'h666;
			{8'd113, 8'd61}: color_data = 12'h666;
			{8'd113, 8'd62}: color_data = 12'h666;
			{8'd113, 8'd63}: color_data = 12'h666;
			{8'd113, 8'd64}: color_data = 12'h666;
			{8'd113, 8'd65}: color_data = 12'h666;
			{8'd113, 8'd66}: color_data = 12'h666;
			{8'd113, 8'd67}: color_data = 12'h666;
			{8'd113, 8'd68}: color_data = 12'h666;
			{8'd113, 8'd69}: color_data = 12'h555;
			{8'd113, 8'd70}: color_data = 12'h555;
			{8'd113, 8'd71}: color_data = 12'h555;
			{8'd113, 8'd72}: color_data = 12'h555;
			{8'd113, 8'd73}: color_data = 12'h555;
			{8'd113, 8'd74}: color_data = 12'h555;
			{8'd113, 8'd75}: color_data = 12'h555;
			{8'd113, 8'd76}: color_data = 12'h555;
			{8'd113, 8'd77}: color_data = 12'h555;
			{8'd113, 8'd78}: color_data = 12'h555;
			{8'd113, 8'd79}: color_data = 12'h555;
			{8'd113, 8'd80}: color_data = 12'h555;
			{8'd113, 8'd81}: color_data = 12'h555;
			{8'd113, 8'd82}: color_data = 12'h444;
			{8'd113, 8'd83}: color_data = 12'h444;
			{8'd113, 8'd84}: color_data = 12'h444;
			{8'd113, 8'd85}: color_data = 12'h444;
			{8'd113, 8'd86}: color_data = 12'h444;
			{8'd113, 8'd87}: color_data = 12'h444;
			{8'd113, 8'd88}: color_data = 12'h444;
			{8'd113, 8'd89}: color_data = 12'h444;
			{8'd113, 8'd90}: color_data = 12'h444;
			{8'd113, 8'd91}: color_data = 12'h444;
			{8'd113, 8'd92}: color_data = 12'h444;
			{8'd113, 8'd93}: color_data = 12'h444;
			{8'd113, 8'd94}: color_data = 12'h444;
			{8'd113, 8'd95}: color_data = 12'h333;
			{8'd113, 8'd96}: color_data = 12'h333;
			{8'd113, 8'd97}: color_data = 12'h333;
			{8'd113, 8'd98}: color_data = 12'h333;
			{8'd113, 8'd99}: color_data = 12'h333;
			{8'd113, 8'd100}: color_data = 12'h333;
			{8'd113, 8'd101}: color_data = 12'h333;
			{8'd113, 8'd102}: color_data = 12'h333;
			{8'd113, 8'd103}: color_data = 12'h333;
			{8'd113, 8'd104}: color_data = 12'h333;
			{8'd113, 8'd105}: color_data = 12'h333;
			{8'd113, 8'd106}: color_data = 12'h333;
			{8'd113, 8'd107}: color_data = 12'h333;
			{8'd113, 8'd108}: color_data = 12'h222;
			{8'd113, 8'd109}: color_data = 12'h222;
			{8'd113, 8'd110}: color_data = 12'h222;
			{8'd113, 8'd111}: color_data = 12'h222;
			{8'd113, 8'd112}: color_data = 12'h222;
			{8'd113, 8'd113}: color_data = 12'h222;
			{8'd113, 8'd114}: color_data = 12'h222;
			{8'd113, 8'd115}: color_data = 12'h222;
			{8'd113, 8'd116}: color_data = 12'h222;
			{8'd113, 8'd117}: color_data = 12'h222;
			{8'd113, 8'd118}: color_data = 12'h222;
			{8'd113, 8'd119}: color_data = 12'h222;
			{8'd113, 8'd120}: color_data = 12'h222;
			{8'd113, 8'd121}: color_data = 12'h222;
			{8'd113, 8'd122}: color_data = 12'h444;
			{8'd113, 8'd123}: color_data = 12'h335;
			{8'd113, 8'd124}: color_data = 12'h34c;
			{8'd113, 8'd125}: color_data = 12'h44d;
			{8'd113, 8'd126}: color_data = 12'h34c;
			{8'd113, 8'd127}: color_data = 12'h779;
			{8'd113, 8'd128}: color_data = 12'haaa;
			{8'd113, 8'd129}: color_data = 12'h888;
			{8'd113, 8'd130}: color_data = 12'h666;
			{8'd113, 8'd131}: color_data = 12'haaa;
			{8'd113, 8'd132}: color_data = 12'hddd;
			{8'd113, 8'd133}: color_data = 12'hfff;
			{8'd113, 8'd134}: color_data = 12'hfff;
			{8'd113, 8'd135}: color_data = 12'hfff;
			{8'd113, 8'd136}: color_data = 12'hfff;
			{8'd113, 8'd137}: color_data = 12'hfff;
			{8'd113, 8'd138}: color_data = 12'hfff;
			{8'd113, 8'd139}: color_data = 12'hfff;
			{8'd113, 8'd140}: color_data = 12'heee;
			{8'd113, 8'd141}: color_data = 12'heee;
			{8'd114, 8'd0}: color_data = 12'hbbb;
			{8'd114, 8'd1}: color_data = 12'hbbb;
			{8'd114, 8'd2}: color_data = 12'hbbb;
			{8'd114, 8'd3}: color_data = 12'hbbb;
			{8'd114, 8'd4}: color_data = 12'haaa;
			{8'd114, 8'd5}: color_data = 12'haaa;
			{8'd114, 8'd6}: color_data = 12'haaa;
			{8'd114, 8'd7}: color_data = 12'haaa;
			{8'd114, 8'd8}: color_data = 12'haaa;
			{8'd114, 8'd9}: color_data = 12'haaa;
			{8'd114, 8'd10}: color_data = 12'haaa;
			{8'd114, 8'd11}: color_data = 12'haaa;
			{8'd114, 8'd12}: color_data = 12'haaa;
			{8'd114, 8'd13}: color_data = 12'haaa;
			{8'd114, 8'd14}: color_data = 12'haaa;
			{8'd114, 8'd15}: color_data = 12'haaa;
			{8'd114, 8'd16}: color_data = 12'h999;
			{8'd114, 8'd17}: color_data = 12'h999;
			{8'd114, 8'd18}: color_data = 12'h999;
			{8'd114, 8'd19}: color_data = 12'h999;
			{8'd114, 8'd20}: color_data = 12'h999;
			{8'd114, 8'd21}: color_data = 12'h999;
			{8'd114, 8'd22}: color_data = 12'h999;
			{8'd114, 8'd23}: color_data = 12'h999;
			{8'd114, 8'd24}: color_data = 12'h999;
			{8'd114, 8'd25}: color_data = 12'h999;
			{8'd114, 8'd26}: color_data = 12'h999;
			{8'd114, 8'd27}: color_data = 12'h999;
			{8'd114, 8'd28}: color_data = 12'h999;
			{8'd114, 8'd29}: color_data = 12'h999;
			{8'd114, 8'd30}: color_data = 12'h999;
			{8'd114, 8'd31}: color_data = 12'h999;
			{8'd114, 8'd32}: color_data = 12'h999;
			{8'd114, 8'd33}: color_data = 12'h888;
			{8'd114, 8'd34}: color_data = 12'h888;
			{8'd114, 8'd35}: color_data = 12'h888;
			{8'd114, 8'd36}: color_data = 12'h888;
			{8'd114, 8'd37}: color_data = 12'h888;
			{8'd114, 8'd38}: color_data = 12'h888;
			{8'd114, 8'd39}: color_data = 12'h888;
			{8'd114, 8'd40}: color_data = 12'h888;
			{8'd114, 8'd41}: color_data = 12'h888;
			{8'd114, 8'd42}: color_data = 12'h888;
			{8'd114, 8'd43}: color_data = 12'h777;
			{8'd114, 8'd44}: color_data = 12'h777;
			{8'd114, 8'd45}: color_data = 12'h777;
			{8'd114, 8'd46}: color_data = 12'h777;
			{8'd114, 8'd47}: color_data = 12'h777;
			{8'd114, 8'd48}: color_data = 12'h777;
			{8'd114, 8'd49}: color_data = 12'h777;
			{8'd114, 8'd50}: color_data = 12'h777;
			{8'd114, 8'd51}: color_data = 12'h777;
			{8'd114, 8'd52}: color_data = 12'h777;
			{8'd114, 8'd53}: color_data = 12'h777;
			{8'd114, 8'd54}: color_data = 12'h777;
			{8'd114, 8'd55}: color_data = 12'h777;
			{8'd114, 8'd56}: color_data = 12'h666;
			{8'd114, 8'd57}: color_data = 12'h666;
			{8'd114, 8'd58}: color_data = 12'h666;
			{8'd114, 8'd59}: color_data = 12'h666;
			{8'd114, 8'd60}: color_data = 12'h666;
			{8'd114, 8'd61}: color_data = 12'h666;
			{8'd114, 8'd62}: color_data = 12'h666;
			{8'd114, 8'd63}: color_data = 12'h666;
			{8'd114, 8'd64}: color_data = 12'h666;
			{8'd114, 8'd65}: color_data = 12'h666;
			{8'd114, 8'd66}: color_data = 12'h666;
			{8'd114, 8'd67}: color_data = 12'h666;
			{8'd114, 8'd68}: color_data = 12'h666;
			{8'd114, 8'd69}: color_data = 12'h555;
			{8'd114, 8'd70}: color_data = 12'h555;
			{8'd114, 8'd71}: color_data = 12'h555;
			{8'd114, 8'd72}: color_data = 12'h555;
			{8'd114, 8'd73}: color_data = 12'h555;
			{8'd114, 8'd74}: color_data = 12'h555;
			{8'd114, 8'd75}: color_data = 12'h555;
			{8'd114, 8'd76}: color_data = 12'h555;
			{8'd114, 8'd77}: color_data = 12'h555;
			{8'd114, 8'd78}: color_data = 12'h555;
			{8'd114, 8'd79}: color_data = 12'h555;
			{8'd114, 8'd80}: color_data = 12'h555;
			{8'd114, 8'd81}: color_data = 12'h555;
			{8'd114, 8'd82}: color_data = 12'h444;
			{8'd114, 8'd83}: color_data = 12'h444;
			{8'd114, 8'd84}: color_data = 12'h444;
			{8'd114, 8'd85}: color_data = 12'h444;
			{8'd114, 8'd86}: color_data = 12'h444;
			{8'd114, 8'd87}: color_data = 12'h444;
			{8'd114, 8'd88}: color_data = 12'h444;
			{8'd114, 8'd89}: color_data = 12'h444;
			{8'd114, 8'd90}: color_data = 12'h444;
			{8'd114, 8'd91}: color_data = 12'h444;
			{8'd114, 8'd92}: color_data = 12'h444;
			{8'd114, 8'd93}: color_data = 12'h444;
			{8'd114, 8'd94}: color_data = 12'h444;
			{8'd114, 8'd95}: color_data = 12'h333;
			{8'd114, 8'd96}: color_data = 12'h333;
			{8'd114, 8'd97}: color_data = 12'h333;
			{8'd114, 8'd98}: color_data = 12'h333;
			{8'd114, 8'd99}: color_data = 12'h333;
			{8'd114, 8'd100}: color_data = 12'h333;
			{8'd114, 8'd101}: color_data = 12'h333;
			{8'd114, 8'd102}: color_data = 12'h333;
			{8'd114, 8'd103}: color_data = 12'h333;
			{8'd114, 8'd104}: color_data = 12'h333;
			{8'd114, 8'd105}: color_data = 12'h333;
			{8'd114, 8'd106}: color_data = 12'h333;
			{8'd114, 8'd107}: color_data = 12'h333;
			{8'd114, 8'd108}: color_data = 12'h333;
			{8'd114, 8'd109}: color_data = 12'h222;
			{8'd114, 8'd110}: color_data = 12'h222;
			{8'd114, 8'd111}: color_data = 12'h222;
			{8'd114, 8'd112}: color_data = 12'h222;
			{8'd114, 8'd113}: color_data = 12'h222;
			{8'd114, 8'd114}: color_data = 12'h222;
			{8'd114, 8'd115}: color_data = 12'h222;
			{8'd114, 8'd116}: color_data = 12'h222;
			{8'd114, 8'd117}: color_data = 12'h222;
			{8'd114, 8'd118}: color_data = 12'h222;
			{8'd114, 8'd119}: color_data = 12'h222;
			{8'd114, 8'd120}: color_data = 12'h222;
			{8'd114, 8'd121}: color_data = 12'h222;
			{8'd114, 8'd122}: color_data = 12'h333;
			{8'd114, 8'd123}: color_data = 12'h348;
			{8'd114, 8'd124}: color_data = 12'h44d;
			{8'd114, 8'd125}: color_data = 12'h34d;
			{8'd114, 8'd126}: color_data = 12'h45a;
			{8'd114, 8'd127}: color_data = 12'h999;
			{8'd114, 8'd128}: color_data = 12'haaa;
			{8'd114, 8'd129}: color_data = 12'h888;
			{8'd114, 8'd130}: color_data = 12'h666;
			{8'd114, 8'd131}: color_data = 12'h999;
			{8'd114, 8'd132}: color_data = 12'hccc;
			{8'd114, 8'd133}: color_data = 12'hfff;
			{8'd114, 8'd134}: color_data = 12'hfff;
			{8'd114, 8'd135}: color_data = 12'hfff;
			{8'd114, 8'd136}: color_data = 12'hfff;
			{8'd114, 8'd137}: color_data = 12'hfff;
			{8'd114, 8'd138}: color_data = 12'hfff;
			{8'd114, 8'd139}: color_data = 12'hfff;
			{8'd114, 8'd140}: color_data = 12'heee;
			{8'd114, 8'd141}: color_data = 12'heee;
			{8'd115, 8'd0}: color_data = 12'hbbb;
			{8'd115, 8'd1}: color_data = 12'hbbb;
			{8'd115, 8'd2}: color_data = 12'hbbb;
			{8'd115, 8'd3}: color_data = 12'hbbb;
			{8'd115, 8'd4}: color_data = 12'haaa;
			{8'd115, 8'd5}: color_data = 12'haaa;
			{8'd115, 8'd6}: color_data = 12'haaa;
			{8'd115, 8'd7}: color_data = 12'haaa;
			{8'd115, 8'd8}: color_data = 12'haaa;
			{8'd115, 8'd9}: color_data = 12'haaa;
			{8'd115, 8'd10}: color_data = 12'haaa;
			{8'd115, 8'd11}: color_data = 12'haaa;
			{8'd115, 8'd12}: color_data = 12'haaa;
			{8'd115, 8'd13}: color_data = 12'haaa;
			{8'd115, 8'd14}: color_data = 12'haaa;
			{8'd115, 8'd15}: color_data = 12'haaa;
			{8'd115, 8'd16}: color_data = 12'h999;
			{8'd115, 8'd17}: color_data = 12'h999;
			{8'd115, 8'd18}: color_data = 12'h999;
			{8'd115, 8'd19}: color_data = 12'h999;
			{8'd115, 8'd20}: color_data = 12'h999;
			{8'd115, 8'd21}: color_data = 12'h999;
			{8'd115, 8'd22}: color_data = 12'h999;
			{8'd115, 8'd23}: color_data = 12'h999;
			{8'd115, 8'd24}: color_data = 12'h999;
			{8'd115, 8'd25}: color_data = 12'h999;
			{8'd115, 8'd26}: color_data = 12'h999;
			{8'd115, 8'd27}: color_data = 12'h999;
			{8'd115, 8'd28}: color_data = 12'h999;
			{8'd115, 8'd29}: color_data = 12'h999;
			{8'd115, 8'd30}: color_data = 12'h888;
			{8'd115, 8'd31}: color_data = 12'h888;
			{8'd115, 8'd32}: color_data = 12'h888;
			{8'd115, 8'd33}: color_data = 12'h888;
			{8'd115, 8'd34}: color_data = 12'h888;
			{8'd115, 8'd35}: color_data = 12'h888;
			{8'd115, 8'd36}: color_data = 12'h888;
			{8'd115, 8'd37}: color_data = 12'h888;
			{8'd115, 8'd38}: color_data = 12'h888;
			{8'd115, 8'd39}: color_data = 12'h888;
			{8'd115, 8'd40}: color_data = 12'h888;
			{8'd115, 8'd41}: color_data = 12'h888;
			{8'd115, 8'd42}: color_data = 12'h888;
			{8'd115, 8'd43}: color_data = 12'h777;
			{8'd115, 8'd44}: color_data = 12'h777;
			{8'd115, 8'd45}: color_data = 12'h777;
			{8'd115, 8'd46}: color_data = 12'h777;
			{8'd115, 8'd47}: color_data = 12'h777;
			{8'd115, 8'd48}: color_data = 12'h777;
			{8'd115, 8'd49}: color_data = 12'h777;
			{8'd115, 8'd50}: color_data = 12'h777;
			{8'd115, 8'd51}: color_data = 12'h777;
			{8'd115, 8'd52}: color_data = 12'h777;
			{8'd115, 8'd53}: color_data = 12'h777;
			{8'd115, 8'd54}: color_data = 12'h777;
			{8'd115, 8'd55}: color_data = 12'h777;
			{8'd115, 8'd56}: color_data = 12'h666;
			{8'd115, 8'd57}: color_data = 12'h666;
			{8'd115, 8'd58}: color_data = 12'h666;
			{8'd115, 8'd59}: color_data = 12'h666;
			{8'd115, 8'd60}: color_data = 12'h666;
			{8'd115, 8'd61}: color_data = 12'h666;
			{8'd115, 8'd62}: color_data = 12'h666;
			{8'd115, 8'd63}: color_data = 12'h666;
			{8'd115, 8'd64}: color_data = 12'h666;
			{8'd115, 8'd65}: color_data = 12'h666;
			{8'd115, 8'd66}: color_data = 12'h666;
			{8'd115, 8'd67}: color_data = 12'h666;
			{8'd115, 8'd68}: color_data = 12'h666;
			{8'd115, 8'd69}: color_data = 12'h555;
			{8'd115, 8'd70}: color_data = 12'h555;
			{8'd115, 8'd71}: color_data = 12'h555;
			{8'd115, 8'd72}: color_data = 12'h555;
			{8'd115, 8'd73}: color_data = 12'h555;
			{8'd115, 8'd74}: color_data = 12'h555;
			{8'd115, 8'd75}: color_data = 12'h555;
			{8'd115, 8'd76}: color_data = 12'h555;
			{8'd115, 8'd77}: color_data = 12'h555;
			{8'd115, 8'd78}: color_data = 12'h555;
			{8'd115, 8'd79}: color_data = 12'h555;
			{8'd115, 8'd80}: color_data = 12'h555;
			{8'd115, 8'd81}: color_data = 12'h555;
			{8'd115, 8'd82}: color_data = 12'h444;
			{8'd115, 8'd83}: color_data = 12'h444;
			{8'd115, 8'd84}: color_data = 12'h444;
			{8'd115, 8'd85}: color_data = 12'h444;
			{8'd115, 8'd86}: color_data = 12'h444;
			{8'd115, 8'd87}: color_data = 12'h444;
			{8'd115, 8'd88}: color_data = 12'h444;
			{8'd115, 8'd89}: color_data = 12'h444;
			{8'd115, 8'd90}: color_data = 12'h444;
			{8'd115, 8'd91}: color_data = 12'h444;
			{8'd115, 8'd92}: color_data = 12'h444;
			{8'd115, 8'd93}: color_data = 12'h444;
			{8'd115, 8'd94}: color_data = 12'h444;
			{8'd115, 8'd95}: color_data = 12'h333;
			{8'd115, 8'd96}: color_data = 12'h333;
			{8'd115, 8'd97}: color_data = 12'h333;
			{8'd115, 8'd98}: color_data = 12'h333;
			{8'd115, 8'd99}: color_data = 12'h333;
			{8'd115, 8'd100}: color_data = 12'h333;
			{8'd115, 8'd101}: color_data = 12'h333;
			{8'd115, 8'd102}: color_data = 12'h333;
			{8'd115, 8'd103}: color_data = 12'h333;
			{8'd115, 8'd104}: color_data = 12'h333;
			{8'd115, 8'd105}: color_data = 12'h333;
			{8'd115, 8'd106}: color_data = 12'h333;
			{8'd115, 8'd107}: color_data = 12'h333;
			{8'd115, 8'd108}: color_data = 12'h333;
			{8'd115, 8'd109}: color_data = 12'h222;
			{8'd115, 8'd110}: color_data = 12'h222;
			{8'd115, 8'd111}: color_data = 12'h222;
			{8'd115, 8'd112}: color_data = 12'h222;
			{8'd115, 8'd113}: color_data = 12'h222;
			{8'd115, 8'd114}: color_data = 12'h222;
			{8'd115, 8'd115}: color_data = 12'h222;
			{8'd115, 8'd116}: color_data = 12'h222;
			{8'd115, 8'd117}: color_data = 12'h222;
			{8'd115, 8'd118}: color_data = 12'h222;
			{8'd115, 8'd119}: color_data = 12'h222;
			{8'd115, 8'd120}: color_data = 12'h222;
			{8'd115, 8'd121}: color_data = 12'h221;
			{8'd115, 8'd122}: color_data = 12'h333;
			{8'd115, 8'd123}: color_data = 12'h449;
			{8'd115, 8'd124}: color_data = 12'h44d;
			{8'd115, 8'd125}: color_data = 12'h34d;
			{8'd115, 8'd126}: color_data = 12'h55a;
			{8'd115, 8'd127}: color_data = 12'haaa;
			{8'd115, 8'd128}: color_data = 12'hbbb;
			{8'd115, 8'd129}: color_data = 12'h999;
			{8'd115, 8'd130}: color_data = 12'h666;
			{8'd115, 8'd131}: color_data = 12'h888;
			{8'd115, 8'd132}: color_data = 12'hccc;
			{8'd115, 8'd133}: color_data = 12'hfff;
			{8'd115, 8'd134}: color_data = 12'hfff;
			{8'd115, 8'd135}: color_data = 12'hfff;
			{8'd115, 8'd136}: color_data = 12'hfff;
			{8'd115, 8'd137}: color_data = 12'hfff;
			{8'd115, 8'd138}: color_data = 12'hfff;
			{8'd115, 8'd139}: color_data = 12'hfff;
			{8'd115, 8'd140}: color_data = 12'hfff;
			{8'd115, 8'd141}: color_data = 12'heee;
			{8'd116, 8'd0}: color_data = 12'hbbb;
			{8'd116, 8'd1}: color_data = 12'hbbb;
			{8'd116, 8'd2}: color_data = 12'hbbb;
			{8'd116, 8'd3}: color_data = 12'hbbb;
			{8'd116, 8'd4}: color_data = 12'haaa;
			{8'd116, 8'd5}: color_data = 12'haaa;
			{8'd116, 8'd6}: color_data = 12'haaa;
			{8'd116, 8'd7}: color_data = 12'haaa;
			{8'd116, 8'd8}: color_data = 12'haaa;
			{8'd116, 8'd9}: color_data = 12'haaa;
			{8'd116, 8'd10}: color_data = 12'haaa;
			{8'd116, 8'd11}: color_data = 12'haaa;
			{8'd116, 8'd12}: color_data = 12'haaa;
			{8'd116, 8'd13}: color_data = 12'haaa;
			{8'd116, 8'd14}: color_data = 12'haaa;
			{8'd116, 8'd15}: color_data = 12'haaa;
			{8'd116, 8'd16}: color_data = 12'h999;
			{8'd116, 8'd17}: color_data = 12'h999;
			{8'd116, 8'd18}: color_data = 12'h999;
			{8'd116, 8'd19}: color_data = 12'h999;
			{8'd116, 8'd20}: color_data = 12'h999;
			{8'd116, 8'd21}: color_data = 12'h999;
			{8'd116, 8'd22}: color_data = 12'h999;
			{8'd116, 8'd23}: color_data = 12'h999;
			{8'd116, 8'd24}: color_data = 12'h999;
			{8'd116, 8'd25}: color_data = 12'h999;
			{8'd116, 8'd26}: color_data = 12'h999;
			{8'd116, 8'd27}: color_data = 12'h999;
			{8'd116, 8'd28}: color_data = 12'h999;
			{8'd116, 8'd29}: color_data = 12'h999;
			{8'd116, 8'd30}: color_data = 12'h888;
			{8'd116, 8'd31}: color_data = 12'h888;
			{8'd116, 8'd32}: color_data = 12'h888;
			{8'd116, 8'd33}: color_data = 12'h888;
			{8'd116, 8'd34}: color_data = 12'h888;
			{8'd116, 8'd35}: color_data = 12'h888;
			{8'd116, 8'd36}: color_data = 12'h888;
			{8'd116, 8'd37}: color_data = 12'h888;
			{8'd116, 8'd38}: color_data = 12'h888;
			{8'd116, 8'd39}: color_data = 12'h888;
			{8'd116, 8'd40}: color_data = 12'h888;
			{8'd116, 8'd41}: color_data = 12'h888;
			{8'd116, 8'd42}: color_data = 12'h888;
			{8'd116, 8'd43}: color_data = 12'h777;
			{8'd116, 8'd44}: color_data = 12'h777;
			{8'd116, 8'd45}: color_data = 12'h777;
			{8'd116, 8'd46}: color_data = 12'h777;
			{8'd116, 8'd47}: color_data = 12'h777;
			{8'd116, 8'd48}: color_data = 12'h777;
			{8'd116, 8'd49}: color_data = 12'h777;
			{8'd116, 8'd50}: color_data = 12'h777;
			{8'd116, 8'd51}: color_data = 12'h777;
			{8'd116, 8'd52}: color_data = 12'h777;
			{8'd116, 8'd53}: color_data = 12'h777;
			{8'd116, 8'd54}: color_data = 12'h777;
			{8'd116, 8'd55}: color_data = 12'h777;
			{8'd116, 8'd56}: color_data = 12'h666;
			{8'd116, 8'd57}: color_data = 12'h666;
			{8'd116, 8'd58}: color_data = 12'h666;
			{8'd116, 8'd59}: color_data = 12'h666;
			{8'd116, 8'd60}: color_data = 12'h666;
			{8'd116, 8'd61}: color_data = 12'h666;
			{8'd116, 8'd62}: color_data = 12'h666;
			{8'd116, 8'd63}: color_data = 12'h666;
			{8'd116, 8'd64}: color_data = 12'h666;
			{8'd116, 8'd65}: color_data = 12'h666;
			{8'd116, 8'd66}: color_data = 12'h666;
			{8'd116, 8'd67}: color_data = 12'h666;
			{8'd116, 8'd68}: color_data = 12'h666;
			{8'd116, 8'd69}: color_data = 12'h555;
			{8'd116, 8'd70}: color_data = 12'h555;
			{8'd116, 8'd71}: color_data = 12'h555;
			{8'd116, 8'd72}: color_data = 12'h555;
			{8'd116, 8'd73}: color_data = 12'h555;
			{8'd116, 8'd74}: color_data = 12'h555;
			{8'd116, 8'd75}: color_data = 12'h555;
			{8'd116, 8'd76}: color_data = 12'h555;
			{8'd116, 8'd77}: color_data = 12'h555;
			{8'd116, 8'd78}: color_data = 12'h555;
			{8'd116, 8'd79}: color_data = 12'h555;
			{8'd116, 8'd80}: color_data = 12'h555;
			{8'd116, 8'd81}: color_data = 12'h555;
			{8'd116, 8'd82}: color_data = 12'h444;
			{8'd116, 8'd83}: color_data = 12'h444;
			{8'd116, 8'd84}: color_data = 12'h444;
			{8'd116, 8'd85}: color_data = 12'h444;
			{8'd116, 8'd86}: color_data = 12'h444;
			{8'd116, 8'd87}: color_data = 12'h444;
			{8'd116, 8'd88}: color_data = 12'h444;
			{8'd116, 8'd89}: color_data = 12'h444;
			{8'd116, 8'd90}: color_data = 12'h444;
			{8'd116, 8'd91}: color_data = 12'h444;
			{8'd116, 8'd92}: color_data = 12'h444;
			{8'd116, 8'd93}: color_data = 12'h444;
			{8'd116, 8'd94}: color_data = 12'h444;
			{8'd116, 8'd95}: color_data = 12'h333;
			{8'd116, 8'd96}: color_data = 12'h333;
			{8'd116, 8'd97}: color_data = 12'h333;
			{8'd116, 8'd98}: color_data = 12'h333;
			{8'd116, 8'd99}: color_data = 12'h333;
			{8'd116, 8'd100}: color_data = 12'h333;
			{8'd116, 8'd101}: color_data = 12'h333;
			{8'd116, 8'd102}: color_data = 12'h333;
			{8'd116, 8'd103}: color_data = 12'h333;
			{8'd116, 8'd104}: color_data = 12'h333;
			{8'd116, 8'd105}: color_data = 12'h333;
			{8'd116, 8'd106}: color_data = 12'h333;
			{8'd116, 8'd107}: color_data = 12'h333;
			{8'd116, 8'd108}: color_data = 12'h333;
			{8'd116, 8'd109}: color_data = 12'h222;
			{8'd116, 8'd110}: color_data = 12'h222;
			{8'd116, 8'd111}: color_data = 12'h222;
			{8'd116, 8'd112}: color_data = 12'h222;
			{8'd116, 8'd113}: color_data = 12'h222;
			{8'd116, 8'd114}: color_data = 12'h222;
			{8'd116, 8'd115}: color_data = 12'h222;
			{8'd116, 8'd116}: color_data = 12'h222;
			{8'd116, 8'd117}: color_data = 12'h222;
			{8'd116, 8'd118}: color_data = 12'h222;
			{8'd116, 8'd119}: color_data = 12'h222;
			{8'd116, 8'd120}: color_data = 12'h222;
			{8'd116, 8'd121}: color_data = 12'h221;
			{8'd116, 8'd122}: color_data = 12'h333;
			{8'd116, 8'd123}: color_data = 12'h349;
			{8'd116, 8'd124}: color_data = 12'h44d;
			{8'd116, 8'd125}: color_data = 12'h44d;
			{8'd116, 8'd126}: color_data = 12'h34c;
			{8'd116, 8'd127}: color_data = 12'h779;
			{8'd116, 8'd128}: color_data = 12'hccc;
			{8'd116, 8'd129}: color_data = 12'h888;
			{8'd116, 8'd130}: color_data = 12'h555;
			{8'd116, 8'd131}: color_data = 12'h888;
			{8'd116, 8'd132}: color_data = 12'hbbb;
			{8'd116, 8'd133}: color_data = 12'hfff;
			{8'd116, 8'd134}: color_data = 12'hfff;
			{8'd116, 8'd135}: color_data = 12'hfff;
			{8'd116, 8'd136}: color_data = 12'hfff;
			{8'd116, 8'd137}: color_data = 12'hfff;
			{8'd116, 8'd138}: color_data = 12'hfff;
			{8'd116, 8'd139}: color_data = 12'hfff;
			{8'd116, 8'd140}: color_data = 12'hfff;
			{8'd116, 8'd141}: color_data = 12'heee;
			{8'd117, 8'd0}: color_data = 12'hbbb;
			{8'd117, 8'd1}: color_data = 12'hbbb;
			{8'd117, 8'd2}: color_data = 12'hbbb;
			{8'd117, 8'd3}: color_data = 12'hbbb;
			{8'd117, 8'd4}: color_data = 12'haaa;
			{8'd117, 8'd5}: color_data = 12'haaa;
			{8'd117, 8'd6}: color_data = 12'haaa;
			{8'd117, 8'd7}: color_data = 12'haaa;
			{8'd117, 8'd8}: color_data = 12'haaa;
			{8'd117, 8'd9}: color_data = 12'haaa;
			{8'd117, 8'd10}: color_data = 12'haaa;
			{8'd117, 8'd11}: color_data = 12'haaa;
			{8'd117, 8'd12}: color_data = 12'haaa;
			{8'd117, 8'd13}: color_data = 12'haaa;
			{8'd117, 8'd14}: color_data = 12'haaa;
			{8'd117, 8'd15}: color_data = 12'haaa;
			{8'd117, 8'd16}: color_data = 12'h999;
			{8'd117, 8'd17}: color_data = 12'h999;
			{8'd117, 8'd18}: color_data = 12'h999;
			{8'd117, 8'd19}: color_data = 12'h999;
			{8'd117, 8'd20}: color_data = 12'h999;
			{8'd117, 8'd21}: color_data = 12'h999;
			{8'd117, 8'd22}: color_data = 12'h999;
			{8'd117, 8'd23}: color_data = 12'h999;
			{8'd117, 8'd24}: color_data = 12'h999;
			{8'd117, 8'd25}: color_data = 12'h999;
			{8'd117, 8'd26}: color_data = 12'h999;
			{8'd117, 8'd27}: color_data = 12'h999;
			{8'd117, 8'd28}: color_data = 12'h999;
			{8'd117, 8'd29}: color_data = 12'h999;
			{8'd117, 8'd30}: color_data = 12'h888;
			{8'd117, 8'd31}: color_data = 12'h888;
			{8'd117, 8'd32}: color_data = 12'h888;
			{8'd117, 8'd33}: color_data = 12'h888;
			{8'd117, 8'd34}: color_data = 12'h888;
			{8'd117, 8'd35}: color_data = 12'h888;
			{8'd117, 8'd36}: color_data = 12'h888;
			{8'd117, 8'd37}: color_data = 12'h888;
			{8'd117, 8'd38}: color_data = 12'h888;
			{8'd117, 8'd39}: color_data = 12'h888;
			{8'd117, 8'd40}: color_data = 12'h888;
			{8'd117, 8'd41}: color_data = 12'h888;
			{8'd117, 8'd42}: color_data = 12'h888;
			{8'd117, 8'd43}: color_data = 12'h777;
			{8'd117, 8'd44}: color_data = 12'h777;
			{8'd117, 8'd45}: color_data = 12'h777;
			{8'd117, 8'd46}: color_data = 12'h777;
			{8'd117, 8'd47}: color_data = 12'h777;
			{8'd117, 8'd48}: color_data = 12'h777;
			{8'd117, 8'd49}: color_data = 12'h777;
			{8'd117, 8'd50}: color_data = 12'h777;
			{8'd117, 8'd51}: color_data = 12'h777;
			{8'd117, 8'd52}: color_data = 12'h777;
			{8'd117, 8'd53}: color_data = 12'h777;
			{8'd117, 8'd54}: color_data = 12'h777;
			{8'd117, 8'd55}: color_data = 12'h777;
			{8'd117, 8'd56}: color_data = 12'h666;
			{8'd117, 8'd57}: color_data = 12'h666;
			{8'd117, 8'd58}: color_data = 12'h666;
			{8'd117, 8'd59}: color_data = 12'h666;
			{8'd117, 8'd60}: color_data = 12'h666;
			{8'd117, 8'd61}: color_data = 12'h666;
			{8'd117, 8'd62}: color_data = 12'h666;
			{8'd117, 8'd63}: color_data = 12'h666;
			{8'd117, 8'd64}: color_data = 12'h666;
			{8'd117, 8'd65}: color_data = 12'h666;
			{8'd117, 8'd66}: color_data = 12'h666;
			{8'd117, 8'd67}: color_data = 12'h666;
			{8'd117, 8'd68}: color_data = 12'h666;
			{8'd117, 8'd69}: color_data = 12'h555;
			{8'd117, 8'd70}: color_data = 12'h555;
			{8'd117, 8'd71}: color_data = 12'h555;
			{8'd117, 8'd72}: color_data = 12'h555;
			{8'd117, 8'd73}: color_data = 12'h555;
			{8'd117, 8'd74}: color_data = 12'h555;
			{8'd117, 8'd75}: color_data = 12'h555;
			{8'd117, 8'd76}: color_data = 12'h555;
			{8'd117, 8'd77}: color_data = 12'h555;
			{8'd117, 8'd78}: color_data = 12'h555;
			{8'd117, 8'd79}: color_data = 12'h555;
			{8'd117, 8'd80}: color_data = 12'h555;
			{8'd117, 8'd81}: color_data = 12'h555;
			{8'd117, 8'd82}: color_data = 12'h444;
			{8'd117, 8'd83}: color_data = 12'h444;
			{8'd117, 8'd84}: color_data = 12'h444;
			{8'd117, 8'd85}: color_data = 12'h444;
			{8'd117, 8'd86}: color_data = 12'h444;
			{8'd117, 8'd87}: color_data = 12'h444;
			{8'd117, 8'd88}: color_data = 12'h444;
			{8'd117, 8'd89}: color_data = 12'h444;
			{8'd117, 8'd90}: color_data = 12'h444;
			{8'd117, 8'd91}: color_data = 12'h444;
			{8'd117, 8'd92}: color_data = 12'h444;
			{8'd117, 8'd93}: color_data = 12'h444;
			{8'd117, 8'd94}: color_data = 12'h444;
			{8'd117, 8'd95}: color_data = 12'h333;
			{8'd117, 8'd96}: color_data = 12'h333;
			{8'd117, 8'd97}: color_data = 12'h333;
			{8'd117, 8'd98}: color_data = 12'h333;
			{8'd117, 8'd99}: color_data = 12'h333;
			{8'd117, 8'd100}: color_data = 12'h333;
			{8'd117, 8'd101}: color_data = 12'h333;
			{8'd117, 8'd102}: color_data = 12'h333;
			{8'd117, 8'd103}: color_data = 12'h333;
			{8'd117, 8'd104}: color_data = 12'h333;
			{8'd117, 8'd105}: color_data = 12'h333;
			{8'd117, 8'd106}: color_data = 12'h333;
			{8'd117, 8'd107}: color_data = 12'h333;
			{8'd117, 8'd108}: color_data = 12'h333;
			{8'd117, 8'd109}: color_data = 12'h222;
			{8'd117, 8'd110}: color_data = 12'h222;
			{8'd117, 8'd111}: color_data = 12'h222;
			{8'd117, 8'd112}: color_data = 12'h222;
			{8'd117, 8'd113}: color_data = 12'h222;
			{8'd117, 8'd114}: color_data = 12'h222;
			{8'd117, 8'd115}: color_data = 12'h222;
			{8'd117, 8'd116}: color_data = 12'h222;
			{8'd117, 8'd117}: color_data = 12'h222;
			{8'd117, 8'd118}: color_data = 12'h222;
			{8'd117, 8'd119}: color_data = 12'h222;
			{8'd117, 8'd120}: color_data = 12'h222;
			{8'd117, 8'd121}: color_data = 12'h222;
			{8'd117, 8'd122}: color_data = 12'h444;
			{8'd117, 8'd123}: color_data = 12'h336;
			{8'd117, 8'd124}: color_data = 12'h44d;
			{8'd117, 8'd125}: color_data = 12'h34d;
			{8'd117, 8'd126}: color_data = 12'h34d;
			{8'd117, 8'd127}: color_data = 12'h44a;
			{8'd117, 8'd128}: color_data = 12'ha89;
			{8'd117, 8'd129}: color_data = 12'h977;
			{8'd117, 8'd130}: color_data = 12'h533;
			{8'd117, 8'd131}: color_data = 12'h888;
			{8'd117, 8'd132}: color_data = 12'hbbb;
			{8'd117, 8'd133}: color_data = 12'heee;
			{8'd117, 8'd134}: color_data = 12'hfff;
			{8'd117, 8'd135}: color_data = 12'hfff;
			{8'd117, 8'd136}: color_data = 12'hfff;
			{8'd117, 8'd137}: color_data = 12'hfff;
			{8'd117, 8'd138}: color_data = 12'hfff;
			{8'd117, 8'd139}: color_data = 12'hfff;
			{8'd117, 8'd140}: color_data = 12'heee;
			{8'd117, 8'd141}: color_data = 12'heee;
			{8'd118, 8'd0}: color_data = 12'hbbb;
			{8'd118, 8'd1}: color_data = 12'hbbb;
			{8'd118, 8'd2}: color_data = 12'hbbb;
			{8'd118, 8'd3}: color_data = 12'hbbb;
			{8'd118, 8'd4}: color_data = 12'haaa;
			{8'd118, 8'd5}: color_data = 12'haaa;
			{8'd118, 8'd6}: color_data = 12'haaa;
			{8'd118, 8'd7}: color_data = 12'haaa;
			{8'd118, 8'd8}: color_data = 12'haaa;
			{8'd118, 8'd9}: color_data = 12'haaa;
			{8'd118, 8'd10}: color_data = 12'haaa;
			{8'd118, 8'd11}: color_data = 12'haaa;
			{8'd118, 8'd12}: color_data = 12'haaa;
			{8'd118, 8'd13}: color_data = 12'haaa;
			{8'd118, 8'd14}: color_data = 12'haaa;
			{8'd118, 8'd15}: color_data = 12'haaa;
			{8'd118, 8'd16}: color_data = 12'h999;
			{8'd118, 8'd17}: color_data = 12'h999;
			{8'd118, 8'd18}: color_data = 12'h999;
			{8'd118, 8'd19}: color_data = 12'h999;
			{8'd118, 8'd20}: color_data = 12'h999;
			{8'd118, 8'd21}: color_data = 12'h999;
			{8'd118, 8'd22}: color_data = 12'h999;
			{8'd118, 8'd23}: color_data = 12'h999;
			{8'd118, 8'd24}: color_data = 12'h999;
			{8'd118, 8'd25}: color_data = 12'h999;
			{8'd118, 8'd26}: color_data = 12'h999;
			{8'd118, 8'd27}: color_data = 12'h999;
			{8'd118, 8'd28}: color_data = 12'h999;
			{8'd118, 8'd29}: color_data = 12'h999;
			{8'd118, 8'd30}: color_data = 12'h888;
			{8'd118, 8'd31}: color_data = 12'h888;
			{8'd118, 8'd32}: color_data = 12'h888;
			{8'd118, 8'd33}: color_data = 12'h888;
			{8'd118, 8'd34}: color_data = 12'h888;
			{8'd118, 8'd35}: color_data = 12'h888;
			{8'd118, 8'd36}: color_data = 12'h888;
			{8'd118, 8'd37}: color_data = 12'h888;
			{8'd118, 8'd38}: color_data = 12'h888;
			{8'd118, 8'd39}: color_data = 12'h888;
			{8'd118, 8'd40}: color_data = 12'h888;
			{8'd118, 8'd41}: color_data = 12'h888;
			{8'd118, 8'd42}: color_data = 12'h888;
			{8'd118, 8'd43}: color_data = 12'h777;
			{8'd118, 8'd44}: color_data = 12'h777;
			{8'd118, 8'd45}: color_data = 12'h777;
			{8'd118, 8'd46}: color_data = 12'h777;
			{8'd118, 8'd47}: color_data = 12'h777;
			{8'd118, 8'd48}: color_data = 12'h777;
			{8'd118, 8'd49}: color_data = 12'h777;
			{8'd118, 8'd50}: color_data = 12'h777;
			{8'd118, 8'd51}: color_data = 12'h777;
			{8'd118, 8'd52}: color_data = 12'h777;
			{8'd118, 8'd53}: color_data = 12'h777;
			{8'd118, 8'd54}: color_data = 12'h777;
			{8'd118, 8'd55}: color_data = 12'h777;
			{8'd118, 8'd56}: color_data = 12'h666;
			{8'd118, 8'd57}: color_data = 12'h666;
			{8'd118, 8'd58}: color_data = 12'h666;
			{8'd118, 8'd59}: color_data = 12'h666;
			{8'd118, 8'd60}: color_data = 12'h666;
			{8'd118, 8'd61}: color_data = 12'h666;
			{8'd118, 8'd62}: color_data = 12'h666;
			{8'd118, 8'd63}: color_data = 12'h666;
			{8'd118, 8'd64}: color_data = 12'h666;
			{8'd118, 8'd65}: color_data = 12'h666;
			{8'd118, 8'd66}: color_data = 12'h666;
			{8'd118, 8'd67}: color_data = 12'h666;
			{8'd118, 8'd68}: color_data = 12'h666;
			{8'd118, 8'd69}: color_data = 12'h555;
			{8'd118, 8'd70}: color_data = 12'h555;
			{8'd118, 8'd71}: color_data = 12'h555;
			{8'd118, 8'd72}: color_data = 12'h555;
			{8'd118, 8'd73}: color_data = 12'h555;
			{8'd118, 8'd74}: color_data = 12'h555;
			{8'd118, 8'd75}: color_data = 12'h555;
			{8'd118, 8'd76}: color_data = 12'h555;
			{8'd118, 8'd77}: color_data = 12'h555;
			{8'd118, 8'd78}: color_data = 12'h555;
			{8'd118, 8'd79}: color_data = 12'h555;
			{8'd118, 8'd80}: color_data = 12'h555;
			{8'd118, 8'd81}: color_data = 12'h555;
			{8'd118, 8'd82}: color_data = 12'h444;
			{8'd118, 8'd83}: color_data = 12'h444;
			{8'd118, 8'd84}: color_data = 12'h444;
			{8'd118, 8'd85}: color_data = 12'h444;
			{8'd118, 8'd86}: color_data = 12'h444;
			{8'd118, 8'd87}: color_data = 12'h444;
			{8'd118, 8'd88}: color_data = 12'h444;
			{8'd118, 8'd89}: color_data = 12'h444;
			{8'd118, 8'd90}: color_data = 12'h444;
			{8'd118, 8'd91}: color_data = 12'h444;
			{8'd118, 8'd92}: color_data = 12'h444;
			{8'd118, 8'd93}: color_data = 12'h444;
			{8'd118, 8'd94}: color_data = 12'h444;
			{8'd118, 8'd95}: color_data = 12'h333;
			{8'd118, 8'd96}: color_data = 12'h333;
			{8'd118, 8'd97}: color_data = 12'h333;
			{8'd118, 8'd98}: color_data = 12'h333;
			{8'd118, 8'd99}: color_data = 12'h333;
			{8'd118, 8'd100}: color_data = 12'h333;
			{8'd118, 8'd101}: color_data = 12'h333;
			{8'd118, 8'd102}: color_data = 12'h333;
			{8'd118, 8'd103}: color_data = 12'h333;
			{8'd118, 8'd104}: color_data = 12'h333;
			{8'd118, 8'd105}: color_data = 12'h333;
			{8'd118, 8'd106}: color_data = 12'h333;
			{8'd118, 8'd107}: color_data = 12'h333;
			{8'd118, 8'd108}: color_data = 12'h333;
			{8'd118, 8'd109}: color_data = 12'h222;
			{8'd118, 8'd110}: color_data = 12'h222;
			{8'd118, 8'd111}: color_data = 12'h222;
			{8'd118, 8'd112}: color_data = 12'h222;
			{8'd118, 8'd113}: color_data = 12'h222;
			{8'd118, 8'd114}: color_data = 12'h222;
			{8'd118, 8'd115}: color_data = 12'h222;
			{8'd118, 8'd116}: color_data = 12'h222;
			{8'd118, 8'd117}: color_data = 12'h222;
			{8'd118, 8'd118}: color_data = 12'h222;
			{8'd118, 8'd119}: color_data = 12'h222;
			{8'd118, 8'd120}: color_data = 12'h222;
			{8'd118, 8'd121}: color_data = 12'h222;
			{8'd118, 8'd122}: color_data = 12'h666;
			{8'd118, 8'd123}: color_data = 12'h556;
			{8'd118, 8'd124}: color_data = 12'h438;
			{8'd118, 8'd125}: color_data = 12'h439;
			{8'd118, 8'd126}: color_data = 12'h646;
			{8'd118, 8'd127}: color_data = 12'h656;
			{8'd118, 8'd128}: color_data = 12'h723;
			{8'd118, 8'd129}: color_data = 12'h812;
			{8'd118, 8'd130}: color_data = 12'h522;
			{8'd118, 8'd131}: color_data = 12'h888;
			{8'd118, 8'd132}: color_data = 12'hbbb;
			{8'd118, 8'd133}: color_data = 12'heee;
			{8'd118, 8'd134}: color_data = 12'hfff;
			{8'd118, 8'd135}: color_data = 12'hfff;
			{8'd118, 8'd136}: color_data = 12'hfff;
			{8'd118, 8'd137}: color_data = 12'hfff;
			{8'd118, 8'd138}: color_data = 12'hfff;
			{8'd118, 8'd139}: color_data = 12'hfff;
			{8'd118, 8'd140}: color_data = 12'heee;
			{8'd118, 8'd141}: color_data = 12'heee;
			{8'd119, 8'd0}: color_data = 12'hbbb;
			{8'd119, 8'd1}: color_data = 12'hbbb;
			{8'd119, 8'd2}: color_data = 12'hbbb;
			{8'd119, 8'd3}: color_data = 12'hbbb;
			{8'd119, 8'd4}: color_data = 12'haaa;
			{8'd119, 8'd5}: color_data = 12'haaa;
			{8'd119, 8'd6}: color_data = 12'haaa;
			{8'd119, 8'd7}: color_data = 12'haaa;
			{8'd119, 8'd8}: color_data = 12'haaa;
			{8'd119, 8'd9}: color_data = 12'haaa;
			{8'd119, 8'd10}: color_data = 12'haaa;
			{8'd119, 8'd11}: color_data = 12'haaa;
			{8'd119, 8'd12}: color_data = 12'haaa;
			{8'd119, 8'd13}: color_data = 12'haaa;
			{8'd119, 8'd14}: color_data = 12'haaa;
			{8'd119, 8'd15}: color_data = 12'haaa;
			{8'd119, 8'd16}: color_data = 12'h999;
			{8'd119, 8'd17}: color_data = 12'h999;
			{8'd119, 8'd18}: color_data = 12'h999;
			{8'd119, 8'd19}: color_data = 12'h999;
			{8'd119, 8'd20}: color_data = 12'h999;
			{8'd119, 8'd21}: color_data = 12'h999;
			{8'd119, 8'd22}: color_data = 12'h999;
			{8'd119, 8'd23}: color_data = 12'h999;
			{8'd119, 8'd24}: color_data = 12'h999;
			{8'd119, 8'd25}: color_data = 12'h999;
			{8'd119, 8'd26}: color_data = 12'h999;
			{8'd119, 8'd27}: color_data = 12'h999;
			{8'd119, 8'd28}: color_data = 12'h999;
			{8'd119, 8'd29}: color_data = 12'h999;
			{8'd119, 8'd30}: color_data = 12'h888;
			{8'd119, 8'd31}: color_data = 12'h888;
			{8'd119, 8'd32}: color_data = 12'h888;
			{8'd119, 8'd33}: color_data = 12'h888;
			{8'd119, 8'd34}: color_data = 12'h888;
			{8'd119, 8'd35}: color_data = 12'h888;
			{8'd119, 8'd36}: color_data = 12'h888;
			{8'd119, 8'd37}: color_data = 12'h888;
			{8'd119, 8'd38}: color_data = 12'h888;
			{8'd119, 8'd39}: color_data = 12'h888;
			{8'd119, 8'd40}: color_data = 12'h888;
			{8'd119, 8'd41}: color_data = 12'h888;
			{8'd119, 8'd42}: color_data = 12'h888;
			{8'd119, 8'd43}: color_data = 12'h777;
			{8'd119, 8'd44}: color_data = 12'h777;
			{8'd119, 8'd45}: color_data = 12'h777;
			{8'd119, 8'd46}: color_data = 12'h777;
			{8'd119, 8'd47}: color_data = 12'h777;
			{8'd119, 8'd48}: color_data = 12'h777;
			{8'd119, 8'd49}: color_data = 12'h777;
			{8'd119, 8'd50}: color_data = 12'h777;
			{8'd119, 8'd51}: color_data = 12'h777;
			{8'd119, 8'd52}: color_data = 12'h777;
			{8'd119, 8'd53}: color_data = 12'h777;
			{8'd119, 8'd54}: color_data = 12'h777;
			{8'd119, 8'd55}: color_data = 12'h777;
			{8'd119, 8'd56}: color_data = 12'h666;
			{8'd119, 8'd57}: color_data = 12'h666;
			{8'd119, 8'd58}: color_data = 12'h666;
			{8'd119, 8'd59}: color_data = 12'h666;
			{8'd119, 8'd60}: color_data = 12'h666;
			{8'd119, 8'd61}: color_data = 12'h666;
			{8'd119, 8'd62}: color_data = 12'h666;
			{8'd119, 8'd63}: color_data = 12'h666;
			{8'd119, 8'd64}: color_data = 12'h666;
			{8'd119, 8'd65}: color_data = 12'h666;
			{8'd119, 8'd66}: color_data = 12'h666;
			{8'd119, 8'd67}: color_data = 12'h666;
			{8'd119, 8'd68}: color_data = 12'h666;
			{8'd119, 8'd69}: color_data = 12'h555;
			{8'd119, 8'd70}: color_data = 12'h555;
			{8'd119, 8'd71}: color_data = 12'h555;
			{8'd119, 8'd72}: color_data = 12'h555;
			{8'd119, 8'd73}: color_data = 12'h555;
			{8'd119, 8'd74}: color_data = 12'h555;
			{8'd119, 8'd75}: color_data = 12'h555;
			{8'd119, 8'd76}: color_data = 12'h555;
			{8'd119, 8'd77}: color_data = 12'h555;
			{8'd119, 8'd78}: color_data = 12'h555;
			{8'd119, 8'd79}: color_data = 12'h555;
			{8'd119, 8'd80}: color_data = 12'h555;
			{8'd119, 8'd81}: color_data = 12'h555;
			{8'd119, 8'd82}: color_data = 12'h444;
			{8'd119, 8'd83}: color_data = 12'h444;
			{8'd119, 8'd84}: color_data = 12'h444;
			{8'd119, 8'd85}: color_data = 12'h444;
			{8'd119, 8'd86}: color_data = 12'h444;
			{8'd119, 8'd87}: color_data = 12'h444;
			{8'd119, 8'd88}: color_data = 12'h444;
			{8'd119, 8'd89}: color_data = 12'h444;
			{8'd119, 8'd90}: color_data = 12'h444;
			{8'd119, 8'd91}: color_data = 12'h444;
			{8'd119, 8'd92}: color_data = 12'h444;
			{8'd119, 8'd93}: color_data = 12'h444;
			{8'd119, 8'd94}: color_data = 12'h444;
			{8'd119, 8'd95}: color_data = 12'h333;
			{8'd119, 8'd96}: color_data = 12'h333;
			{8'd119, 8'd97}: color_data = 12'h333;
			{8'd119, 8'd98}: color_data = 12'h333;
			{8'd119, 8'd99}: color_data = 12'h333;
			{8'd119, 8'd100}: color_data = 12'h333;
			{8'd119, 8'd101}: color_data = 12'h333;
			{8'd119, 8'd102}: color_data = 12'h333;
			{8'd119, 8'd103}: color_data = 12'h333;
			{8'd119, 8'd104}: color_data = 12'h333;
			{8'd119, 8'd105}: color_data = 12'h333;
			{8'd119, 8'd106}: color_data = 12'h333;
			{8'd119, 8'd107}: color_data = 12'h333;
			{8'd119, 8'd108}: color_data = 12'h333;
			{8'd119, 8'd109}: color_data = 12'h222;
			{8'd119, 8'd110}: color_data = 12'h222;
			{8'd119, 8'd111}: color_data = 12'h222;
			{8'd119, 8'd112}: color_data = 12'h222;
			{8'd119, 8'd113}: color_data = 12'h222;
			{8'd119, 8'd114}: color_data = 12'h222;
			{8'd119, 8'd115}: color_data = 12'h222;
			{8'd119, 8'd116}: color_data = 12'h222;
			{8'd119, 8'd117}: color_data = 12'h222;
			{8'd119, 8'd118}: color_data = 12'h222;
			{8'd119, 8'd119}: color_data = 12'h222;
			{8'd119, 8'd120}: color_data = 12'h222;
			{8'd119, 8'd121}: color_data = 12'h222;
			{8'd119, 8'd122}: color_data = 12'h665;
			{8'd119, 8'd123}: color_data = 12'h755;
			{8'd119, 8'd124}: color_data = 12'h722;
			{8'd119, 8'd125}: color_data = 12'h733;
			{8'd119, 8'd126}: color_data = 12'ha75;
			{8'd119, 8'd127}: color_data = 12'hb85;
			{8'd119, 8'd128}: color_data = 12'h964;
			{8'd119, 8'd129}: color_data = 12'h712;
			{8'd119, 8'd130}: color_data = 12'h422;
			{8'd119, 8'd131}: color_data = 12'h888;
			{8'd119, 8'd132}: color_data = 12'hbbb;
			{8'd119, 8'd133}: color_data = 12'heee;
			{8'd119, 8'd134}: color_data = 12'hfff;
			{8'd119, 8'd135}: color_data = 12'hfff;
			{8'd119, 8'd136}: color_data = 12'hfff;
			{8'd119, 8'd137}: color_data = 12'hfff;
			{8'd119, 8'd138}: color_data = 12'hfff;
			{8'd119, 8'd139}: color_data = 12'hfff;
			{8'd119, 8'd140}: color_data = 12'heee;
			{8'd119, 8'd141}: color_data = 12'heee;
			{8'd120, 8'd0}: color_data = 12'hbbb;
			{8'd120, 8'd1}: color_data = 12'hbbb;
			{8'd120, 8'd2}: color_data = 12'hbbb;
			{8'd120, 8'd3}: color_data = 12'hbbb;
			{8'd120, 8'd4}: color_data = 12'haaa;
			{8'd120, 8'd5}: color_data = 12'haaa;
			{8'd120, 8'd6}: color_data = 12'haaa;
			{8'd120, 8'd7}: color_data = 12'haaa;
			{8'd120, 8'd8}: color_data = 12'haaa;
			{8'd120, 8'd9}: color_data = 12'haaa;
			{8'd120, 8'd10}: color_data = 12'haaa;
			{8'd120, 8'd11}: color_data = 12'haaa;
			{8'd120, 8'd12}: color_data = 12'haaa;
			{8'd120, 8'd13}: color_data = 12'haaa;
			{8'd120, 8'd14}: color_data = 12'haaa;
			{8'd120, 8'd15}: color_data = 12'haaa;
			{8'd120, 8'd16}: color_data = 12'h999;
			{8'd120, 8'd17}: color_data = 12'h999;
			{8'd120, 8'd18}: color_data = 12'h999;
			{8'd120, 8'd19}: color_data = 12'h999;
			{8'd120, 8'd20}: color_data = 12'h999;
			{8'd120, 8'd21}: color_data = 12'h999;
			{8'd120, 8'd22}: color_data = 12'h999;
			{8'd120, 8'd23}: color_data = 12'h999;
			{8'd120, 8'd24}: color_data = 12'h999;
			{8'd120, 8'd25}: color_data = 12'h999;
			{8'd120, 8'd26}: color_data = 12'h999;
			{8'd120, 8'd27}: color_data = 12'h999;
			{8'd120, 8'd28}: color_data = 12'h999;
			{8'd120, 8'd29}: color_data = 12'h999;
			{8'd120, 8'd30}: color_data = 12'h888;
			{8'd120, 8'd31}: color_data = 12'h888;
			{8'd120, 8'd32}: color_data = 12'h888;
			{8'd120, 8'd33}: color_data = 12'h888;
			{8'd120, 8'd34}: color_data = 12'h888;
			{8'd120, 8'd35}: color_data = 12'h888;
			{8'd120, 8'd36}: color_data = 12'h888;
			{8'd120, 8'd37}: color_data = 12'h888;
			{8'd120, 8'd38}: color_data = 12'h888;
			{8'd120, 8'd39}: color_data = 12'h888;
			{8'd120, 8'd40}: color_data = 12'h888;
			{8'd120, 8'd41}: color_data = 12'h888;
			{8'd120, 8'd42}: color_data = 12'h888;
			{8'd120, 8'd43}: color_data = 12'h777;
			{8'd120, 8'd44}: color_data = 12'h777;
			{8'd120, 8'd45}: color_data = 12'h777;
			{8'd120, 8'd46}: color_data = 12'h777;
			{8'd120, 8'd47}: color_data = 12'h777;
			{8'd120, 8'd48}: color_data = 12'h777;
			{8'd120, 8'd49}: color_data = 12'h777;
			{8'd120, 8'd50}: color_data = 12'h777;
			{8'd120, 8'd51}: color_data = 12'h777;
			{8'd120, 8'd52}: color_data = 12'h777;
			{8'd120, 8'd53}: color_data = 12'h777;
			{8'd120, 8'd54}: color_data = 12'h777;
			{8'd120, 8'd55}: color_data = 12'h777;
			{8'd120, 8'd56}: color_data = 12'h666;
			{8'd120, 8'd57}: color_data = 12'h666;
			{8'd120, 8'd58}: color_data = 12'h666;
			{8'd120, 8'd59}: color_data = 12'h666;
			{8'd120, 8'd60}: color_data = 12'h666;
			{8'd120, 8'd61}: color_data = 12'h666;
			{8'd120, 8'd62}: color_data = 12'h666;
			{8'd120, 8'd63}: color_data = 12'h666;
			{8'd120, 8'd64}: color_data = 12'h666;
			{8'd120, 8'd65}: color_data = 12'h666;
			{8'd120, 8'd66}: color_data = 12'h666;
			{8'd120, 8'd67}: color_data = 12'h666;
			{8'd120, 8'd68}: color_data = 12'h666;
			{8'd120, 8'd69}: color_data = 12'h555;
			{8'd120, 8'd70}: color_data = 12'h555;
			{8'd120, 8'd71}: color_data = 12'h555;
			{8'd120, 8'd72}: color_data = 12'h555;
			{8'd120, 8'd73}: color_data = 12'h555;
			{8'd120, 8'd74}: color_data = 12'h555;
			{8'd120, 8'd75}: color_data = 12'h555;
			{8'd120, 8'd76}: color_data = 12'h555;
			{8'd120, 8'd77}: color_data = 12'h555;
			{8'd120, 8'd78}: color_data = 12'h555;
			{8'd120, 8'd79}: color_data = 12'h555;
			{8'd120, 8'd80}: color_data = 12'h555;
			{8'd120, 8'd81}: color_data = 12'h555;
			{8'd120, 8'd82}: color_data = 12'h444;
			{8'd120, 8'd83}: color_data = 12'h444;
			{8'd120, 8'd84}: color_data = 12'h444;
			{8'd120, 8'd85}: color_data = 12'h444;
			{8'd120, 8'd86}: color_data = 12'h444;
			{8'd120, 8'd87}: color_data = 12'h444;
			{8'd120, 8'd88}: color_data = 12'h444;
			{8'd120, 8'd89}: color_data = 12'h444;
			{8'd120, 8'd90}: color_data = 12'h444;
			{8'd120, 8'd91}: color_data = 12'h444;
			{8'd120, 8'd92}: color_data = 12'h444;
			{8'd120, 8'd93}: color_data = 12'h444;
			{8'd120, 8'd94}: color_data = 12'h444;
			{8'd120, 8'd95}: color_data = 12'h333;
			{8'd120, 8'd96}: color_data = 12'h333;
			{8'd120, 8'd97}: color_data = 12'h333;
			{8'd120, 8'd98}: color_data = 12'h333;
			{8'd120, 8'd99}: color_data = 12'h333;
			{8'd120, 8'd100}: color_data = 12'h333;
			{8'd120, 8'd101}: color_data = 12'h333;
			{8'd120, 8'd102}: color_data = 12'h333;
			{8'd120, 8'd103}: color_data = 12'h333;
			{8'd120, 8'd104}: color_data = 12'h333;
			{8'd120, 8'd105}: color_data = 12'h333;
			{8'd120, 8'd106}: color_data = 12'h333;
			{8'd120, 8'd107}: color_data = 12'h333;
			{8'd120, 8'd108}: color_data = 12'h333;
			{8'd120, 8'd109}: color_data = 12'h222;
			{8'd120, 8'd110}: color_data = 12'h222;
			{8'd120, 8'd111}: color_data = 12'h222;
			{8'd120, 8'd112}: color_data = 12'h222;
			{8'd120, 8'd113}: color_data = 12'h222;
			{8'd120, 8'd114}: color_data = 12'h222;
			{8'd120, 8'd115}: color_data = 12'h222;
			{8'd120, 8'd116}: color_data = 12'h222;
			{8'd120, 8'd117}: color_data = 12'h222;
			{8'd120, 8'd118}: color_data = 12'h222;
			{8'd120, 8'd119}: color_data = 12'h222;
			{8'd120, 8'd120}: color_data = 12'h222;
			{8'd120, 8'd121}: color_data = 12'h222;
			{8'd120, 8'd122}: color_data = 12'h432;
			{8'd120, 8'd123}: color_data = 12'h822;
			{8'd120, 8'd124}: color_data = 12'hb23;
			{8'd120, 8'd125}: color_data = 12'h843;
			{8'd120, 8'd126}: color_data = 12'hb86;
			{8'd120, 8'd127}: color_data = 12'hb75;
			{8'd120, 8'd128}: color_data = 12'hb85;
			{8'd120, 8'd129}: color_data = 12'h522;
			{8'd120, 8'd130}: color_data = 12'h322;
			{8'd120, 8'd131}: color_data = 12'h888;
			{8'd120, 8'd132}: color_data = 12'hbbb;
			{8'd120, 8'd133}: color_data = 12'hfff;
			{8'd120, 8'd134}: color_data = 12'hfff;
			{8'd120, 8'd135}: color_data = 12'hfff;
			{8'd120, 8'd136}: color_data = 12'hfff;
			{8'd120, 8'd137}: color_data = 12'hfff;
			{8'd120, 8'd138}: color_data = 12'hfff;
			{8'd120, 8'd139}: color_data = 12'hfff;
			{8'd120, 8'd140}: color_data = 12'heee;
			{8'd120, 8'd141}: color_data = 12'hddd;
			{8'd121, 8'd0}: color_data = 12'hbbb;
			{8'd121, 8'd1}: color_data = 12'hbbb;
			{8'd121, 8'd2}: color_data = 12'hbbb;
			{8'd121, 8'd3}: color_data = 12'hbbb;
			{8'd121, 8'd4}: color_data = 12'haaa;
			{8'd121, 8'd5}: color_data = 12'haaa;
			{8'd121, 8'd6}: color_data = 12'haaa;
			{8'd121, 8'd7}: color_data = 12'haaa;
			{8'd121, 8'd8}: color_data = 12'haaa;
			{8'd121, 8'd9}: color_data = 12'haaa;
			{8'd121, 8'd10}: color_data = 12'haaa;
			{8'd121, 8'd11}: color_data = 12'haaa;
			{8'd121, 8'd12}: color_data = 12'haaa;
			{8'd121, 8'd13}: color_data = 12'haaa;
			{8'd121, 8'd14}: color_data = 12'haaa;
			{8'd121, 8'd15}: color_data = 12'haaa;
			{8'd121, 8'd16}: color_data = 12'h999;
			{8'd121, 8'd17}: color_data = 12'h999;
			{8'd121, 8'd18}: color_data = 12'h999;
			{8'd121, 8'd19}: color_data = 12'h999;
			{8'd121, 8'd20}: color_data = 12'h999;
			{8'd121, 8'd21}: color_data = 12'h999;
			{8'd121, 8'd22}: color_data = 12'h999;
			{8'd121, 8'd23}: color_data = 12'h999;
			{8'd121, 8'd24}: color_data = 12'h999;
			{8'd121, 8'd25}: color_data = 12'h999;
			{8'd121, 8'd26}: color_data = 12'h999;
			{8'd121, 8'd27}: color_data = 12'h999;
			{8'd121, 8'd28}: color_data = 12'h999;
			{8'd121, 8'd29}: color_data = 12'h999;
			{8'd121, 8'd30}: color_data = 12'h888;
			{8'd121, 8'd31}: color_data = 12'h888;
			{8'd121, 8'd32}: color_data = 12'h888;
			{8'd121, 8'd33}: color_data = 12'h888;
			{8'd121, 8'd34}: color_data = 12'h888;
			{8'd121, 8'd35}: color_data = 12'h888;
			{8'd121, 8'd36}: color_data = 12'h888;
			{8'd121, 8'd37}: color_data = 12'h888;
			{8'd121, 8'd38}: color_data = 12'h888;
			{8'd121, 8'd39}: color_data = 12'h888;
			{8'd121, 8'd40}: color_data = 12'h888;
			{8'd121, 8'd41}: color_data = 12'h888;
			{8'd121, 8'd42}: color_data = 12'h888;
			{8'd121, 8'd43}: color_data = 12'h777;
			{8'd121, 8'd44}: color_data = 12'h777;
			{8'd121, 8'd45}: color_data = 12'h777;
			{8'd121, 8'd46}: color_data = 12'h777;
			{8'd121, 8'd47}: color_data = 12'h777;
			{8'd121, 8'd48}: color_data = 12'h777;
			{8'd121, 8'd49}: color_data = 12'h777;
			{8'd121, 8'd50}: color_data = 12'h777;
			{8'd121, 8'd51}: color_data = 12'h777;
			{8'd121, 8'd52}: color_data = 12'h777;
			{8'd121, 8'd53}: color_data = 12'h777;
			{8'd121, 8'd54}: color_data = 12'h777;
			{8'd121, 8'd55}: color_data = 12'h777;
			{8'd121, 8'd56}: color_data = 12'h666;
			{8'd121, 8'd57}: color_data = 12'h666;
			{8'd121, 8'd58}: color_data = 12'h666;
			{8'd121, 8'd59}: color_data = 12'h666;
			{8'd121, 8'd60}: color_data = 12'h666;
			{8'd121, 8'd61}: color_data = 12'h666;
			{8'd121, 8'd62}: color_data = 12'h666;
			{8'd121, 8'd63}: color_data = 12'h666;
			{8'd121, 8'd64}: color_data = 12'h666;
			{8'd121, 8'd65}: color_data = 12'h666;
			{8'd121, 8'd66}: color_data = 12'h666;
			{8'd121, 8'd67}: color_data = 12'h666;
			{8'd121, 8'd68}: color_data = 12'h666;
			{8'd121, 8'd69}: color_data = 12'h555;
			{8'd121, 8'd70}: color_data = 12'h555;
			{8'd121, 8'd71}: color_data = 12'h555;
			{8'd121, 8'd72}: color_data = 12'h555;
			{8'd121, 8'd73}: color_data = 12'h555;
			{8'd121, 8'd74}: color_data = 12'h555;
			{8'd121, 8'd75}: color_data = 12'h555;
			{8'd121, 8'd76}: color_data = 12'h555;
			{8'd121, 8'd77}: color_data = 12'h555;
			{8'd121, 8'd78}: color_data = 12'h555;
			{8'd121, 8'd79}: color_data = 12'h555;
			{8'd121, 8'd80}: color_data = 12'h555;
			{8'd121, 8'd81}: color_data = 12'h555;
			{8'd121, 8'd82}: color_data = 12'h444;
			{8'd121, 8'd83}: color_data = 12'h444;
			{8'd121, 8'd84}: color_data = 12'h444;
			{8'd121, 8'd85}: color_data = 12'h444;
			{8'd121, 8'd86}: color_data = 12'h444;
			{8'd121, 8'd87}: color_data = 12'h444;
			{8'd121, 8'd88}: color_data = 12'h444;
			{8'd121, 8'd89}: color_data = 12'h444;
			{8'd121, 8'd90}: color_data = 12'h444;
			{8'd121, 8'd91}: color_data = 12'h444;
			{8'd121, 8'd92}: color_data = 12'h444;
			{8'd121, 8'd93}: color_data = 12'h444;
			{8'd121, 8'd94}: color_data = 12'h444;
			{8'd121, 8'd95}: color_data = 12'h333;
			{8'd121, 8'd96}: color_data = 12'h333;
			{8'd121, 8'd97}: color_data = 12'h333;
			{8'd121, 8'd98}: color_data = 12'h333;
			{8'd121, 8'd99}: color_data = 12'h333;
			{8'd121, 8'd100}: color_data = 12'h333;
			{8'd121, 8'd101}: color_data = 12'h333;
			{8'd121, 8'd102}: color_data = 12'h333;
			{8'd121, 8'd103}: color_data = 12'h333;
			{8'd121, 8'd104}: color_data = 12'h333;
			{8'd121, 8'd105}: color_data = 12'h333;
			{8'd121, 8'd106}: color_data = 12'h333;
			{8'd121, 8'd107}: color_data = 12'h333;
			{8'd121, 8'd108}: color_data = 12'h333;
			{8'd121, 8'd109}: color_data = 12'h222;
			{8'd121, 8'd110}: color_data = 12'h222;
			{8'd121, 8'd111}: color_data = 12'h222;
			{8'd121, 8'd112}: color_data = 12'h222;
			{8'd121, 8'd113}: color_data = 12'h222;
			{8'd121, 8'd114}: color_data = 12'h222;
			{8'd121, 8'd115}: color_data = 12'h222;
			{8'd121, 8'd116}: color_data = 12'h222;
			{8'd121, 8'd117}: color_data = 12'h222;
			{8'd121, 8'd118}: color_data = 12'h222;
			{8'd121, 8'd119}: color_data = 12'h222;
			{8'd121, 8'd120}: color_data = 12'h222;
			{8'd121, 8'd121}: color_data = 12'h122;
			{8'd121, 8'd122}: color_data = 12'h422;
			{8'd121, 8'd123}: color_data = 12'h822;
			{8'd121, 8'd124}: color_data = 12'ha23;
			{8'd121, 8'd125}: color_data = 12'h733;
			{8'd121, 8'd126}: color_data = 12'h974;
			{8'd121, 8'd127}: color_data = 12'hb85;
			{8'd121, 8'd128}: color_data = 12'hc96;
			{8'd121, 8'd129}: color_data = 12'h753;
			{8'd121, 8'd130}: color_data = 12'h322;
			{8'd121, 8'd131}: color_data = 12'h999;
			{8'd121, 8'd132}: color_data = 12'hccc;
			{8'd121, 8'd133}: color_data = 12'hfff;
			{8'd121, 8'd134}: color_data = 12'hfff;
			{8'd121, 8'd135}: color_data = 12'hfff;
			{8'd121, 8'd136}: color_data = 12'hfff;
			{8'd121, 8'd137}: color_data = 12'hfff;
			{8'd121, 8'd138}: color_data = 12'hfff;
			{8'd121, 8'd139}: color_data = 12'hfff;
			{8'd121, 8'd140}: color_data = 12'heee;
			{8'd121, 8'd141}: color_data = 12'hddd;
			{8'd122, 8'd0}: color_data = 12'hbbb;
			{8'd122, 8'd1}: color_data = 12'hbbb;
			{8'd122, 8'd2}: color_data = 12'hbbb;
			{8'd122, 8'd3}: color_data = 12'hbbb;
			{8'd122, 8'd4}: color_data = 12'haaa;
			{8'd122, 8'd5}: color_data = 12'haaa;
			{8'd122, 8'd6}: color_data = 12'haaa;
			{8'd122, 8'd7}: color_data = 12'haaa;
			{8'd122, 8'd8}: color_data = 12'haaa;
			{8'd122, 8'd9}: color_data = 12'haaa;
			{8'd122, 8'd10}: color_data = 12'haaa;
			{8'd122, 8'd11}: color_data = 12'haaa;
			{8'd122, 8'd12}: color_data = 12'haaa;
			{8'd122, 8'd13}: color_data = 12'haaa;
			{8'd122, 8'd14}: color_data = 12'haaa;
			{8'd122, 8'd15}: color_data = 12'haaa;
			{8'd122, 8'd16}: color_data = 12'h999;
			{8'd122, 8'd17}: color_data = 12'h999;
			{8'd122, 8'd18}: color_data = 12'h999;
			{8'd122, 8'd19}: color_data = 12'h999;
			{8'd122, 8'd20}: color_data = 12'h999;
			{8'd122, 8'd21}: color_data = 12'h999;
			{8'd122, 8'd22}: color_data = 12'h999;
			{8'd122, 8'd23}: color_data = 12'h999;
			{8'd122, 8'd24}: color_data = 12'h999;
			{8'd122, 8'd25}: color_data = 12'h999;
			{8'd122, 8'd26}: color_data = 12'h999;
			{8'd122, 8'd27}: color_data = 12'h999;
			{8'd122, 8'd28}: color_data = 12'h999;
			{8'd122, 8'd29}: color_data = 12'h999;
			{8'd122, 8'd30}: color_data = 12'h888;
			{8'd122, 8'd31}: color_data = 12'h888;
			{8'd122, 8'd32}: color_data = 12'h888;
			{8'd122, 8'd33}: color_data = 12'h888;
			{8'd122, 8'd34}: color_data = 12'h888;
			{8'd122, 8'd35}: color_data = 12'h888;
			{8'd122, 8'd36}: color_data = 12'h888;
			{8'd122, 8'd37}: color_data = 12'h888;
			{8'd122, 8'd38}: color_data = 12'h888;
			{8'd122, 8'd39}: color_data = 12'h888;
			{8'd122, 8'd40}: color_data = 12'h888;
			{8'd122, 8'd41}: color_data = 12'h888;
			{8'd122, 8'd42}: color_data = 12'h888;
			{8'd122, 8'd43}: color_data = 12'h777;
			{8'd122, 8'd44}: color_data = 12'h777;
			{8'd122, 8'd45}: color_data = 12'h777;
			{8'd122, 8'd46}: color_data = 12'h777;
			{8'd122, 8'd47}: color_data = 12'h777;
			{8'd122, 8'd48}: color_data = 12'h777;
			{8'd122, 8'd49}: color_data = 12'h777;
			{8'd122, 8'd50}: color_data = 12'h777;
			{8'd122, 8'd51}: color_data = 12'h777;
			{8'd122, 8'd52}: color_data = 12'h777;
			{8'd122, 8'd53}: color_data = 12'h777;
			{8'd122, 8'd54}: color_data = 12'h777;
			{8'd122, 8'd55}: color_data = 12'h777;
			{8'd122, 8'd56}: color_data = 12'h666;
			{8'd122, 8'd57}: color_data = 12'h666;
			{8'd122, 8'd58}: color_data = 12'h666;
			{8'd122, 8'd59}: color_data = 12'h666;
			{8'd122, 8'd60}: color_data = 12'h666;
			{8'd122, 8'd61}: color_data = 12'h666;
			{8'd122, 8'd62}: color_data = 12'h666;
			{8'd122, 8'd63}: color_data = 12'h666;
			{8'd122, 8'd64}: color_data = 12'h666;
			{8'd122, 8'd65}: color_data = 12'h666;
			{8'd122, 8'd66}: color_data = 12'h666;
			{8'd122, 8'd67}: color_data = 12'h666;
			{8'd122, 8'd68}: color_data = 12'h666;
			{8'd122, 8'd69}: color_data = 12'h555;
			{8'd122, 8'd70}: color_data = 12'h555;
			{8'd122, 8'd71}: color_data = 12'h555;
			{8'd122, 8'd72}: color_data = 12'h555;
			{8'd122, 8'd73}: color_data = 12'h555;
			{8'd122, 8'd74}: color_data = 12'h555;
			{8'd122, 8'd75}: color_data = 12'h555;
			{8'd122, 8'd76}: color_data = 12'h555;
			{8'd122, 8'd77}: color_data = 12'h555;
			{8'd122, 8'd78}: color_data = 12'h555;
			{8'd122, 8'd79}: color_data = 12'h555;
			{8'd122, 8'd80}: color_data = 12'h555;
			{8'd122, 8'd81}: color_data = 12'h555;
			{8'd122, 8'd82}: color_data = 12'h444;
			{8'd122, 8'd83}: color_data = 12'h444;
			{8'd122, 8'd84}: color_data = 12'h444;
			{8'd122, 8'd85}: color_data = 12'h444;
			{8'd122, 8'd86}: color_data = 12'h444;
			{8'd122, 8'd87}: color_data = 12'h444;
			{8'd122, 8'd88}: color_data = 12'h444;
			{8'd122, 8'd89}: color_data = 12'h444;
			{8'd122, 8'd90}: color_data = 12'h444;
			{8'd122, 8'd91}: color_data = 12'h444;
			{8'd122, 8'd92}: color_data = 12'h444;
			{8'd122, 8'd93}: color_data = 12'h444;
			{8'd122, 8'd94}: color_data = 12'h444;
			{8'd122, 8'd95}: color_data = 12'h333;
			{8'd122, 8'd96}: color_data = 12'h333;
			{8'd122, 8'd97}: color_data = 12'h333;
			{8'd122, 8'd98}: color_data = 12'h333;
			{8'd122, 8'd99}: color_data = 12'h333;
			{8'd122, 8'd100}: color_data = 12'h333;
			{8'd122, 8'd101}: color_data = 12'h333;
			{8'd122, 8'd102}: color_data = 12'h333;
			{8'd122, 8'd103}: color_data = 12'h333;
			{8'd122, 8'd104}: color_data = 12'h333;
			{8'd122, 8'd105}: color_data = 12'h333;
			{8'd122, 8'd106}: color_data = 12'h333;
			{8'd122, 8'd107}: color_data = 12'h333;
			{8'd122, 8'd108}: color_data = 12'h333;
			{8'd122, 8'd109}: color_data = 12'h222;
			{8'd122, 8'd110}: color_data = 12'h222;
			{8'd122, 8'd111}: color_data = 12'h222;
			{8'd122, 8'd112}: color_data = 12'h222;
			{8'd122, 8'd113}: color_data = 12'h222;
			{8'd122, 8'd114}: color_data = 12'h222;
			{8'd122, 8'd115}: color_data = 12'h222;
			{8'd122, 8'd116}: color_data = 12'h222;
			{8'd122, 8'd117}: color_data = 12'h222;
			{8'd122, 8'd118}: color_data = 12'h222;
			{8'd122, 8'd119}: color_data = 12'h222;
			{8'd122, 8'd120}: color_data = 12'h122;
			{8'd122, 8'd121}: color_data = 12'h222;
			{8'd122, 8'd122}: color_data = 12'h622;
			{8'd122, 8'd123}: color_data = 12'h922;
			{8'd122, 8'd124}: color_data = 12'hb33;
			{8'd122, 8'd125}: color_data = 12'h733;
			{8'd122, 8'd126}: color_data = 12'h532;
			{8'd122, 8'd127}: color_data = 12'h753;
			{8'd122, 8'd128}: color_data = 12'hc96;
			{8'd122, 8'd129}: color_data = 12'ha75;
			{8'd122, 8'd130}: color_data = 12'h433;
			{8'd122, 8'd131}: color_data = 12'h999;
			{8'd122, 8'd132}: color_data = 12'hccc;
			{8'd122, 8'd133}: color_data = 12'hfff;
			{8'd122, 8'd134}: color_data = 12'hfff;
			{8'd122, 8'd135}: color_data = 12'hfff;
			{8'd122, 8'd136}: color_data = 12'hfff;
			{8'd122, 8'd137}: color_data = 12'hfff;
			{8'd122, 8'd138}: color_data = 12'hfff;
			{8'd122, 8'd139}: color_data = 12'hfff;
			{8'd122, 8'd140}: color_data = 12'hddd;
			{8'd122, 8'd141}: color_data = 12'hddd;
			{8'd123, 8'd0}: color_data = 12'hbbb;
			{8'd123, 8'd1}: color_data = 12'hbbb;
			{8'd123, 8'd2}: color_data = 12'hbbb;
			{8'd123, 8'd3}: color_data = 12'hbbb;
			{8'd123, 8'd4}: color_data = 12'haaa;
			{8'd123, 8'd5}: color_data = 12'haaa;
			{8'd123, 8'd6}: color_data = 12'haaa;
			{8'd123, 8'd7}: color_data = 12'haaa;
			{8'd123, 8'd8}: color_data = 12'haaa;
			{8'd123, 8'd9}: color_data = 12'haaa;
			{8'd123, 8'd10}: color_data = 12'haaa;
			{8'd123, 8'd11}: color_data = 12'haaa;
			{8'd123, 8'd12}: color_data = 12'haaa;
			{8'd123, 8'd13}: color_data = 12'haaa;
			{8'd123, 8'd14}: color_data = 12'haaa;
			{8'd123, 8'd15}: color_data = 12'haaa;
			{8'd123, 8'd16}: color_data = 12'h999;
			{8'd123, 8'd17}: color_data = 12'h999;
			{8'd123, 8'd18}: color_data = 12'h999;
			{8'd123, 8'd19}: color_data = 12'h999;
			{8'd123, 8'd20}: color_data = 12'h999;
			{8'd123, 8'd21}: color_data = 12'h999;
			{8'd123, 8'd22}: color_data = 12'h999;
			{8'd123, 8'd23}: color_data = 12'h999;
			{8'd123, 8'd24}: color_data = 12'h999;
			{8'd123, 8'd25}: color_data = 12'h999;
			{8'd123, 8'd26}: color_data = 12'h999;
			{8'd123, 8'd27}: color_data = 12'h999;
			{8'd123, 8'd28}: color_data = 12'h999;
			{8'd123, 8'd29}: color_data = 12'h999;
			{8'd123, 8'd30}: color_data = 12'h888;
			{8'd123, 8'd31}: color_data = 12'h888;
			{8'd123, 8'd32}: color_data = 12'h888;
			{8'd123, 8'd33}: color_data = 12'h888;
			{8'd123, 8'd34}: color_data = 12'h888;
			{8'd123, 8'd35}: color_data = 12'h888;
			{8'd123, 8'd36}: color_data = 12'h888;
			{8'd123, 8'd37}: color_data = 12'h888;
			{8'd123, 8'd38}: color_data = 12'h888;
			{8'd123, 8'd39}: color_data = 12'h888;
			{8'd123, 8'd40}: color_data = 12'h888;
			{8'd123, 8'd41}: color_data = 12'h888;
			{8'd123, 8'd42}: color_data = 12'h888;
			{8'd123, 8'd43}: color_data = 12'h777;
			{8'd123, 8'd44}: color_data = 12'h777;
			{8'd123, 8'd45}: color_data = 12'h777;
			{8'd123, 8'd46}: color_data = 12'h777;
			{8'd123, 8'd47}: color_data = 12'h777;
			{8'd123, 8'd48}: color_data = 12'h777;
			{8'd123, 8'd49}: color_data = 12'h777;
			{8'd123, 8'd50}: color_data = 12'h777;
			{8'd123, 8'd51}: color_data = 12'h777;
			{8'd123, 8'd52}: color_data = 12'h777;
			{8'd123, 8'd53}: color_data = 12'h777;
			{8'd123, 8'd54}: color_data = 12'h777;
			{8'd123, 8'd55}: color_data = 12'h777;
			{8'd123, 8'd56}: color_data = 12'h666;
			{8'd123, 8'd57}: color_data = 12'h666;
			{8'd123, 8'd58}: color_data = 12'h666;
			{8'd123, 8'd59}: color_data = 12'h666;
			{8'd123, 8'd60}: color_data = 12'h666;
			{8'd123, 8'd61}: color_data = 12'h666;
			{8'd123, 8'd62}: color_data = 12'h666;
			{8'd123, 8'd63}: color_data = 12'h666;
			{8'd123, 8'd64}: color_data = 12'h666;
			{8'd123, 8'd65}: color_data = 12'h666;
			{8'd123, 8'd66}: color_data = 12'h666;
			{8'd123, 8'd67}: color_data = 12'h666;
			{8'd123, 8'd68}: color_data = 12'h666;
			{8'd123, 8'd69}: color_data = 12'h555;
			{8'd123, 8'd70}: color_data = 12'h555;
			{8'd123, 8'd71}: color_data = 12'h555;
			{8'd123, 8'd72}: color_data = 12'h555;
			{8'd123, 8'd73}: color_data = 12'h555;
			{8'd123, 8'd74}: color_data = 12'h555;
			{8'd123, 8'd75}: color_data = 12'h555;
			{8'd123, 8'd76}: color_data = 12'h555;
			{8'd123, 8'd77}: color_data = 12'h555;
			{8'd123, 8'd78}: color_data = 12'h555;
			{8'd123, 8'd79}: color_data = 12'h555;
			{8'd123, 8'd80}: color_data = 12'h555;
			{8'd123, 8'd81}: color_data = 12'h555;
			{8'd123, 8'd82}: color_data = 12'h444;
			{8'd123, 8'd83}: color_data = 12'h444;
			{8'd123, 8'd84}: color_data = 12'h444;
			{8'd123, 8'd85}: color_data = 12'h444;
			{8'd123, 8'd86}: color_data = 12'h444;
			{8'd123, 8'd87}: color_data = 12'h444;
			{8'd123, 8'd88}: color_data = 12'h444;
			{8'd123, 8'd89}: color_data = 12'h444;
			{8'd123, 8'd90}: color_data = 12'h444;
			{8'd123, 8'd91}: color_data = 12'h444;
			{8'd123, 8'd92}: color_data = 12'h444;
			{8'd123, 8'd93}: color_data = 12'h444;
			{8'd123, 8'd94}: color_data = 12'h444;
			{8'd123, 8'd95}: color_data = 12'h333;
			{8'd123, 8'd96}: color_data = 12'h333;
			{8'd123, 8'd97}: color_data = 12'h333;
			{8'd123, 8'd98}: color_data = 12'h333;
			{8'd123, 8'd99}: color_data = 12'h333;
			{8'd123, 8'd100}: color_data = 12'h333;
			{8'd123, 8'd101}: color_data = 12'h333;
			{8'd123, 8'd102}: color_data = 12'h333;
			{8'd123, 8'd103}: color_data = 12'h333;
			{8'd123, 8'd104}: color_data = 12'h333;
			{8'd123, 8'd105}: color_data = 12'h333;
			{8'd123, 8'd106}: color_data = 12'h333;
			{8'd123, 8'd107}: color_data = 12'h333;
			{8'd123, 8'd108}: color_data = 12'h333;
			{8'd123, 8'd109}: color_data = 12'h222;
			{8'd123, 8'd110}: color_data = 12'h222;
			{8'd123, 8'd111}: color_data = 12'h222;
			{8'd123, 8'd112}: color_data = 12'h222;
			{8'd123, 8'd113}: color_data = 12'h222;
			{8'd123, 8'd114}: color_data = 12'h222;
			{8'd123, 8'd115}: color_data = 12'h222;
			{8'd123, 8'd116}: color_data = 12'h222;
			{8'd123, 8'd117}: color_data = 12'h222;
			{8'd123, 8'd118}: color_data = 12'h222;
			{8'd123, 8'd119}: color_data = 12'h222;
			{8'd123, 8'd120}: color_data = 12'h222;
			{8'd123, 8'd121}: color_data = 12'h522;
			{8'd123, 8'd122}: color_data = 12'h923;
			{8'd123, 8'd123}: color_data = 12'hb34;
			{8'd123, 8'd124}: color_data = 12'hb34;
			{8'd123, 8'd125}: color_data = 12'h833;
			{8'd123, 8'd126}: color_data = 12'h864;
			{8'd123, 8'd127}: color_data = 12'ha75;
			{8'd123, 8'd128}: color_data = 12'h975;
			{8'd123, 8'd129}: color_data = 12'h754;
			{8'd123, 8'd130}: color_data = 12'h754;
			{8'd123, 8'd131}: color_data = 12'haaa;
			{8'd123, 8'd132}: color_data = 12'hddd;
			{8'd123, 8'd133}: color_data = 12'hfff;
			{8'd123, 8'd134}: color_data = 12'hfff;
			{8'd123, 8'd135}: color_data = 12'hfff;
			{8'd123, 8'd136}: color_data = 12'hfff;
			{8'd123, 8'd137}: color_data = 12'hfff;
			{8'd123, 8'd138}: color_data = 12'hfff;
			{8'd123, 8'd139}: color_data = 12'hfff;
			{8'd123, 8'd140}: color_data = 12'hddd;
			{8'd123, 8'd141}: color_data = 12'hccc;
			{8'd124, 8'd0}: color_data = 12'hbbb;
			{8'd124, 8'd1}: color_data = 12'hbbb;
			{8'd124, 8'd2}: color_data = 12'hbbb;
			{8'd124, 8'd3}: color_data = 12'hbbb;
			{8'd124, 8'd4}: color_data = 12'haaa;
			{8'd124, 8'd5}: color_data = 12'haaa;
			{8'd124, 8'd6}: color_data = 12'haaa;
			{8'd124, 8'd7}: color_data = 12'haaa;
			{8'd124, 8'd8}: color_data = 12'haaa;
			{8'd124, 8'd9}: color_data = 12'haaa;
			{8'd124, 8'd10}: color_data = 12'haaa;
			{8'd124, 8'd11}: color_data = 12'haaa;
			{8'd124, 8'd12}: color_data = 12'haaa;
			{8'd124, 8'd13}: color_data = 12'haaa;
			{8'd124, 8'd14}: color_data = 12'haaa;
			{8'd124, 8'd15}: color_data = 12'haaa;
			{8'd124, 8'd16}: color_data = 12'h999;
			{8'd124, 8'd17}: color_data = 12'h999;
			{8'd124, 8'd18}: color_data = 12'h999;
			{8'd124, 8'd19}: color_data = 12'h999;
			{8'd124, 8'd20}: color_data = 12'h999;
			{8'd124, 8'd21}: color_data = 12'h999;
			{8'd124, 8'd22}: color_data = 12'h999;
			{8'd124, 8'd23}: color_data = 12'h999;
			{8'd124, 8'd24}: color_data = 12'h999;
			{8'd124, 8'd25}: color_data = 12'h999;
			{8'd124, 8'd26}: color_data = 12'h999;
			{8'd124, 8'd27}: color_data = 12'h999;
			{8'd124, 8'd28}: color_data = 12'h999;
			{8'd124, 8'd29}: color_data = 12'h999;
			{8'd124, 8'd30}: color_data = 12'h888;
			{8'd124, 8'd31}: color_data = 12'h888;
			{8'd124, 8'd32}: color_data = 12'h888;
			{8'd124, 8'd33}: color_data = 12'h888;
			{8'd124, 8'd34}: color_data = 12'h888;
			{8'd124, 8'd35}: color_data = 12'h888;
			{8'd124, 8'd36}: color_data = 12'h888;
			{8'd124, 8'd37}: color_data = 12'h888;
			{8'd124, 8'd38}: color_data = 12'h888;
			{8'd124, 8'd39}: color_data = 12'h888;
			{8'd124, 8'd40}: color_data = 12'h888;
			{8'd124, 8'd41}: color_data = 12'h888;
			{8'd124, 8'd42}: color_data = 12'h888;
			{8'd124, 8'd43}: color_data = 12'h777;
			{8'd124, 8'd44}: color_data = 12'h777;
			{8'd124, 8'd45}: color_data = 12'h777;
			{8'd124, 8'd46}: color_data = 12'h777;
			{8'd124, 8'd47}: color_data = 12'h777;
			{8'd124, 8'd48}: color_data = 12'h777;
			{8'd124, 8'd49}: color_data = 12'h777;
			{8'd124, 8'd50}: color_data = 12'h777;
			{8'd124, 8'd51}: color_data = 12'h777;
			{8'd124, 8'd52}: color_data = 12'h777;
			{8'd124, 8'd53}: color_data = 12'h777;
			{8'd124, 8'd54}: color_data = 12'h777;
			{8'd124, 8'd55}: color_data = 12'h777;
			{8'd124, 8'd56}: color_data = 12'h666;
			{8'd124, 8'd57}: color_data = 12'h666;
			{8'd124, 8'd58}: color_data = 12'h666;
			{8'd124, 8'd59}: color_data = 12'h666;
			{8'd124, 8'd60}: color_data = 12'h666;
			{8'd124, 8'd61}: color_data = 12'h666;
			{8'd124, 8'd62}: color_data = 12'h666;
			{8'd124, 8'd63}: color_data = 12'h666;
			{8'd124, 8'd64}: color_data = 12'h666;
			{8'd124, 8'd65}: color_data = 12'h666;
			{8'd124, 8'd66}: color_data = 12'h666;
			{8'd124, 8'd67}: color_data = 12'h666;
			{8'd124, 8'd68}: color_data = 12'h666;
			{8'd124, 8'd69}: color_data = 12'h555;
			{8'd124, 8'd70}: color_data = 12'h555;
			{8'd124, 8'd71}: color_data = 12'h555;
			{8'd124, 8'd72}: color_data = 12'h555;
			{8'd124, 8'd73}: color_data = 12'h555;
			{8'd124, 8'd74}: color_data = 12'h555;
			{8'd124, 8'd75}: color_data = 12'h555;
			{8'd124, 8'd76}: color_data = 12'h555;
			{8'd124, 8'd77}: color_data = 12'h555;
			{8'd124, 8'd78}: color_data = 12'h555;
			{8'd124, 8'd79}: color_data = 12'h555;
			{8'd124, 8'd80}: color_data = 12'h555;
			{8'd124, 8'd81}: color_data = 12'h555;
			{8'd124, 8'd82}: color_data = 12'h444;
			{8'd124, 8'd83}: color_data = 12'h444;
			{8'd124, 8'd84}: color_data = 12'h444;
			{8'd124, 8'd85}: color_data = 12'h444;
			{8'd124, 8'd86}: color_data = 12'h444;
			{8'd124, 8'd87}: color_data = 12'h444;
			{8'd124, 8'd88}: color_data = 12'h444;
			{8'd124, 8'd89}: color_data = 12'h444;
			{8'd124, 8'd90}: color_data = 12'h444;
			{8'd124, 8'd91}: color_data = 12'h444;
			{8'd124, 8'd92}: color_data = 12'h444;
			{8'd124, 8'd93}: color_data = 12'h444;
			{8'd124, 8'd94}: color_data = 12'h444;
			{8'd124, 8'd95}: color_data = 12'h333;
			{8'd124, 8'd96}: color_data = 12'h333;
			{8'd124, 8'd97}: color_data = 12'h333;
			{8'd124, 8'd98}: color_data = 12'h333;
			{8'd124, 8'd99}: color_data = 12'h333;
			{8'd124, 8'd100}: color_data = 12'h333;
			{8'd124, 8'd101}: color_data = 12'h333;
			{8'd124, 8'd102}: color_data = 12'h333;
			{8'd124, 8'd103}: color_data = 12'h333;
			{8'd124, 8'd104}: color_data = 12'h333;
			{8'd124, 8'd105}: color_data = 12'h333;
			{8'd124, 8'd106}: color_data = 12'h333;
			{8'd124, 8'd107}: color_data = 12'h333;
			{8'd124, 8'd108}: color_data = 12'h333;
			{8'd124, 8'd109}: color_data = 12'h222;
			{8'd124, 8'd110}: color_data = 12'h222;
			{8'd124, 8'd111}: color_data = 12'h222;
			{8'd124, 8'd112}: color_data = 12'h222;
			{8'd124, 8'd113}: color_data = 12'h222;
			{8'd124, 8'd114}: color_data = 12'h222;
			{8'd124, 8'd115}: color_data = 12'h222;
			{8'd124, 8'd116}: color_data = 12'h222;
			{8'd124, 8'd117}: color_data = 12'h222;
			{8'd124, 8'd118}: color_data = 12'h222;
			{8'd124, 8'd119}: color_data = 12'h222;
			{8'd124, 8'd120}: color_data = 12'h622;
			{8'd124, 8'd121}: color_data = 12'h923;
			{8'd124, 8'd122}: color_data = 12'hb34;
			{8'd124, 8'd123}: color_data = 12'hb34;
			{8'd124, 8'd124}: color_data = 12'ha23;
			{8'd124, 8'd125}: color_data = 12'h733;
			{8'd124, 8'd126}: color_data = 12'ha85;
			{8'd124, 8'd127}: color_data = 12'hb86;
			{8'd124, 8'd128}: color_data = 12'h433;
			{8'd124, 8'd129}: color_data = 12'h221;
			{8'd124, 8'd130}: color_data = 12'h544;
			{8'd124, 8'd131}: color_data = 12'hbbb;
			{8'd124, 8'd132}: color_data = 12'heee;
			{8'd124, 8'd133}: color_data = 12'hfff;
			{8'd124, 8'd134}: color_data = 12'hfff;
			{8'd124, 8'd135}: color_data = 12'hfff;
			{8'd124, 8'd136}: color_data = 12'hfff;
			{8'd124, 8'd137}: color_data = 12'hfff;
			{8'd124, 8'd138}: color_data = 12'hfff;
			{8'd124, 8'd139}: color_data = 12'hfff;
			{8'd124, 8'd140}: color_data = 12'hccc;
			{8'd124, 8'd141}: color_data = 12'hbbb;
			{8'd125, 8'd0}: color_data = 12'hbbb;
			{8'd125, 8'd1}: color_data = 12'hbbb;
			{8'd125, 8'd2}: color_data = 12'hbbb;
			{8'd125, 8'd3}: color_data = 12'hbbb;
			{8'd125, 8'd4}: color_data = 12'haaa;
			{8'd125, 8'd5}: color_data = 12'haaa;
			{8'd125, 8'd6}: color_data = 12'haaa;
			{8'd125, 8'd7}: color_data = 12'haaa;
			{8'd125, 8'd8}: color_data = 12'haaa;
			{8'd125, 8'd9}: color_data = 12'haaa;
			{8'd125, 8'd10}: color_data = 12'haaa;
			{8'd125, 8'd11}: color_data = 12'haaa;
			{8'd125, 8'd12}: color_data = 12'haaa;
			{8'd125, 8'd13}: color_data = 12'haaa;
			{8'd125, 8'd14}: color_data = 12'haaa;
			{8'd125, 8'd15}: color_data = 12'haaa;
			{8'd125, 8'd16}: color_data = 12'h999;
			{8'd125, 8'd17}: color_data = 12'h999;
			{8'd125, 8'd18}: color_data = 12'h999;
			{8'd125, 8'd19}: color_data = 12'h999;
			{8'd125, 8'd20}: color_data = 12'h999;
			{8'd125, 8'd21}: color_data = 12'h999;
			{8'd125, 8'd22}: color_data = 12'h999;
			{8'd125, 8'd23}: color_data = 12'h999;
			{8'd125, 8'd24}: color_data = 12'h999;
			{8'd125, 8'd25}: color_data = 12'h999;
			{8'd125, 8'd26}: color_data = 12'h999;
			{8'd125, 8'd27}: color_data = 12'h999;
			{8'd125, 8'd28}: color_data = 12'h999;
			{8'd125, 8'd29}: color_data = 12'h999;
			{8'd125, 8'd30}: color_data = 12'h888;
			{8'd125, 8'd31}: color_data = 12'h888;
			{8'd125, 8'd32}: color_data = 12'h888;
			{8'd125, 8'd33}: color_data = 12'h888;
			{8'd125, 8'd34}: color_data = 12'h888;
			{8'd125, 8'd35}: color_data = 12'h888;
			{8'd125, 8'd36}: color_data = 12'h888;
			{8'd125, 8'd37}: color_data = 12'h888;
			{8'd125, 8'd38}: color_data = 12'h888;
			{8'd125, 8'd39}: color_data = 12'h888;
			{8'd125, 8'd40}: color_data = 12'h888;
			{8'd125, 8'd41}: color_data = 12'h888;
			{8'd125, 8'd42}: color_data = 12'h888;
			{8'd125, 8'd43}: color_data = 12'h777;
			{8'd125, 8'd44}: color_data = 12'h777;
			{8'd125, 8'd45}: color_data = 12'h777;
			{8'd125, 8'd46}: color_data = 12'h777;
			{8'd125, 8'd47}: color_data = 12'h777;
			{8'd125, 8'd48}: color_data = 12'h777;
			{8'd125, 8'd49}: color_data = 12'h777;
			{8'd125, 8'd50}: color_data = 12'h777;
			{8'd125, 8'd51}: color_data = 12'h777;
			{8'd125, 8'd52}: color_data = 12'h777;
			{8'd125, 8'd53}: color_data = 12'h777;
			{8'd125, 8'd54}: color_data = 12'h777;
			{8'd125, 8'd55}: color_data = 12'h777;
			{8'd125, 8'd56}: color_data = 12'h666;
			{8'd125, 8'd57}: color_data = 12'h666;
			{8'd125, 8'd58}: color_data = 12'h666;
			{8'd125, 8'd59}: color_data = 12'h666;
			{8'd125, 8'd60}: color_data = 12'h666;
			{8'd125, 8'd61}: color_data = 12'h666;
			{8'd125, 8'd62}: color_data = 12'h666;
			{8'd125, 8'd63}: color_data = 12'h666;
			{8'd125, 8'd64}: color_data = 12'h666;
			{8'd125, 8'd65}: color_data = 12'h666;
			{8'd125, 8'd66}: color_data = 12'h666;
			{8'd125, 8'd67}: color_data = 12'h666;
			{8'd125, 8'd68}: color_data = 12'h666;
			{8'd125, 8'd69}: color_data = 12'h555;
			{8'd125, 8'd70}: color_data = 12'h555;
			{8'd125, 8'd71}: color_data = 12'h555;
			{8'd125, 8'd72}: color_data = 12'h555;
			{8'd125, 8'd73}: color_data = 12'h555;
			{8'd125, 8'd74}: color_data = 12'h555;
			{8'd125, 8'd75}: color_data = 12'h555;
			{8'd125, 8'd76}: color_data = 12'h555;
			{8'd125, 8'd77}: color_data = 12'h555;
			{8'd125, 8'd78}: color_data = 12'h555;
			{8'd125, 8'd79}: color_data = 12'h555;
			{8'd125, 8'd80}: color_data = 12'h555;
			{8'd125, 8'd81}: color_data = 12'h555;
			{8'd125, 8'd82}: color_data = 12'h444;
			{8'd125, 8'd83}: color_data = 12'h444;
			{8'd125, 8'd84}: color_data = 12'h444;
			{8'd125, 8'd85}: color_data = 12'h444;
			{8'd125, 8'd86}: color_data = 12'h444;
			{8'd125, 8'd87}: color_data = 12'h444;
			{8'd125, 8'd88}: color_data = 12'h444;
			{8'd125, 8'd89}: color_data = 12'h444;
			{8'd125, 8'd90}: color_data = 12'h444;
			{8'd125, 8'd91}: color_data = 12'h444;
			{8'd125, 8'd92}: color_data = 12'h444;
			{8'd125, 8'd93}: color_data = 12'h444;
			{8'd125, 8'd94}: color_data = 12'h444;
			{8'd125, 8'd95}: color_data = 12'h333;
			{8'd125, 8'd96}: color_data = 12'h333;
			{8'd125, 8'd97}: color_data = 12'h333;
			{8'd125, 8'd98}: color_data = 12'h333;
			{8'd125, 8'd99}: color_data = 12'h333;
			{8'd125, 8'd100}: color_data = 12'h333;
			{8'd125, 8'd101}: color_data = 12'h333;
			{8'd125, 8'd102}: color_data = 12'h333;
			{8'd125, 8'd103}: color_data = 12'h333;
			{8'd125, 8'd104}: color_data = 12'h333;
			{8'd125, 8'd105}: color_data = 12'h333;
			{8'd125, 8'd106}: color_data = 12'h333;
			{8'd125, 8'd107}: color_data = 12'h333;
			{8'd125, 8'd108}: color_data = 12'h333;
			{8'd125, 8'd109}: color_data = 12'h222;
			{8'd125, 8'd110}: color_data = 12'h222;
			{8'd125, 8'd111}: color_data = 12'h222;
			{8'd125, 8'd112}: color_data = 12'h222;
			{8'd125, 8'd113}: color_data = 12'h222;
			{8'd125, 8'd114}: color_data = 12'h222;
			{8'd125, 8'd115}: color_data = 12'h222;
			{8'd125, 8'd116}: color_data = 12'h222;
			{8'd125, 8'd117}: color_data = 12'h222;
			{8'd125, 8'd118}: color_data = 12'h222;
			{8'd125, 8'd119}: color_data = 12'h422;
			{8'd125, 8'd120}: color_data = 12'h822;
			{8'd125, 8'd121}: color_data = 12'hb34;
			{8'd125, 8'd122}: color_data = 12'hb34;
			{8'd125, 8'd123}: color_data = 12'hb23;
			{8'd125, 8'd124}: color_data = 12'ha23;
			{8'd125, 8'd125}: color_data = 12'h533;
			{8'd125, 8'd126}: color_data = 12'h653;
			{8'd125, 8'd127}: color_data = 12'h974;
			{8'd125, 8'd128}: color_data = 12'h865;
			{8'd125, 8'd129}: color_data = 12'h221;
			{8'd125, 8'd130}: color_data = 12'h433;
			{8'd125, 8'd131}: color_data = 12'hccc;
			{8'd125, 8'd132}: color_data = 12'heee;
			{8'd125, 8'd133}: color_data = 12'hfff;
			{8'd125, 8'd134}: color_data = 12'hfff;
			{8'd125, 8'd135}: color_data = 12'hfff;
			{8'd125, 8'd136}: color_data = 12'hfff;
			{8'd125, 8'd137}: color_data = 12'hfff;
			{8'd125, 8'd138}: color_data = 12'hfff;
			{8'd125, 8'd139}: color_data = 12'hfff;
			{8'd125, 8'd140}: color_data = 12'hccc;
			{8'd125, 8'd141}: color_data = 12'h999;
			{8'd126, 8'd0}: color_data = 12'hbbb;
			{8'd126, 8'd1}: color_data = 12'hbbb;
			{8'd126, 8'd2}: color_data = 12'hbbb;
			{8'd126, 8'd3}: color_data = 12'hbbb;
			{8'd126, 8'd4}: color_data = 12'haaa;
			{8'd126, 8'd5}: color_data = 12'haaa;
			{8'd126, 8'd6}: color_data = 12'haaa;
			{8'd126, 8'd7}: color_data = 12'haaa;
			{8'd126, 8'd8}: color_data = 12'haaa;
			{8'd126, 8'd9}: color_data = 12'haaa;
			{8'd126, 8'd10}: color_data = 12'haaa;
			{8'd126, 8'd11}: color_data = 12'haaa;
			{8'd126, 8'd12}: color_data = 12'haaa;
			{8'd126, 8'd13}: color_data = 12'haaa;
			{8'd126, 8'd14}: color_data = 12'haaa;
			{8'd126, 8'd15}: color_data = 12'haaa;
			{8'd126, 8'd16}: color_data = 12'haaa;
			{8'd126, 8'd17}: color_data = 12'h999;
			{8'd126, 8'd18}: color_data = 12'h999;
			{8'd126, 8'd19}: color_data = 12'h999;
			{8'd126, 8'd20}: color_data = 12'h999;
			{8'd126, 8'd21}: color_data = 12'h999;
			{8'd126, 8'd22}: color_data = 12'h999;
			{8'd126, 8'd23}: color_data = 12'h999;
			{8'd126, 8'd24}: color_data = 12'h999;
			{8'd126, 8'd25}: color_data = 12'h999;
			{8'd126, 8'd26}: color_data = 12'h999;
			{8'd126, 8'd27}: color_data = 12'h999;
			{8'd126, 8'd28}: color_data = 12'h999;
			{8'd126, 8'd29}: color_data = 12'h999;
			{8'd126, 8'd30}: color_data = 12'h888;
			{8'd126, 8'd31}: color_data = 12'h888;
			{8'd126, 8'd32}: color_data = 12'h888;
			{8'd126, 8'd33}: color_data = 12'h888;
			{8'd126, 8'd34}: color_data = 12'h888;
			{8'd126, 8'd35}: color_data = 12'h888;
			{8'd126, 8'd36}: color_data = 12'h888;
			{8'd126, 8'd37}: color_data = 12'h888;
			{8'd126, 8'd38}: color_data = 12'h888;
			{8'd126, 8'd39}: color_data = 12'h888;
			{8'd126, 8'd40}: color_data = 12'h888;
			{8'd126, 8'd41}: color_data = 12'h888;
			{8'd126, 8'd42}: color_data = 12'h888;
			{8'd126, 8'd43}: color_data = 12'h888;
			{8'd126, 8'd44}: color_data = 12'h777;
			{8'd126, 8'd45}: color_data = 12'h777;
			{8'd126, 8'd46}: color_data = 12'h777;
			{8'd126, 8'd47}: color_data = 12'h777;
			{8'd126, 8'd48}: color_data = 12'h777;
			{8'd126, 8'd49}: color_data = 12'h777;
			{8'd126, 8'd50}: color_data = 12'h777;
			{8'd126, 8'd51}: color_data = 12'h777;
			{8'd126, 8'd52}: color_data = 12'h777;
			{8'd126, 8'd53}: color_data = 12'h777;
			{8'd126, 8'd54}: color_data = 12'h777;
			{8'd126, 8'd55}: color_data = 12'h777;
			{8'd126, 8'd56}: color_data = 12'h666;
			{8'd126, 8'd57}: color_data = 12'h666;
			{8'd126, 8'd58}: color_data = 12'h666;
			{8'd126, 8'd59}: color_data = 12'h666;
			{8'd126, 8'd60}: color_data = 12'h666;
			{8'd126, 8'd61}: color_data = 12'h666;
			{8'd126, 8'd62}: color_data = 12'h666;
			{8'd126, 8'd63}: color_data = 12'h666;
			{8'd126, 8'd64}: color_data = 12'h666;
			{8'd126, 8'd65}: color_data = 12'h666;
			{8'd126, 8'd66}: color_data = 12'h666;
			{8'd126, 8'd67}: color_data = 12'h666;
			{8'd126, 8'd68}: color_data = 12'h666;
			{8'd126, 8'd69}: color_data = 12'h555;
			{8'd126, 8'd70}: color_data = 12'h555;
			{8'd126, 8'd71}: color_data = 12'h555;
			{8'd126, 8'd72}: color_data = 12'h555;
			{8'd126, 8'd73}: color_data = 12'h555;
			{8'd126, 8'd74}: color_data = 12'h555;
			{8'd126, 8'd75}: color_data = 12'h555;
			{8'd126, 8'd76}: color_data = 12'h555;
			{8'd126, 8'd77}: color_data = 12'h555;
			{8'd126, 8'd78}: color_data = 12'h555;
			{8'd126, 8'd79}: color_data = 12'h555;
			{8'd126, 8'd80}: color_data = 12'h555;
			{8'd126, 8'd81}: color_data = 12'h555;
			{8'd126, 8'd82}: color_data = 12'h444;
			{8'd126, 8'd83}: color_data = 12'h444;
			{8'd126, 8'd84}: color_data = 12'h444;
			{8'd126, 8'd85}: color_data = 12'h444;
			{8'd126, 8'd86}: color_data = 12'h444;
			{8'd126, 8'd87}: color_data = 12'h444;
			{8'd126, 8'd88}: color_data = 12'h444;
			{8'd126, 8'd89}: color_data = 12'h444;
			{8'd126, 8'd90}: color_data = 12'h444;
			{8'd126, 8'd91}: color_data = 12'h444;
			{8'd126, 8'd92}: color_data = 12'h444;
			{8'd126, 8'd93}: color_data = 12'h444;
			{8'd126, 8'd94}: color_data = 12'h444;
			{8'd126, 8'd95}: color_data = 12'h333;
			{8'd126, 8'd96}: color_data = 12'h333;
			{8'd126, 8'd97}: color_data = 12'h333;
			{8'd126, 8'd98}: color_data = 12'h333;
			{8'd126, 8'd99}: color_data = 12'h333;
			{8'd126, 8'd100}: color_data = 12'h333;
			{8'd126, 8'd101}: color_data = 12'h333;
			{8'd126, 8'd102}: color_data = 12'h333;
			{8'd126, 8'd103}: color_data = 12'h333;
			{8'd126, 8'd104}: color_data = 12'h333;
			{8'd126, 8'd105}: color_data = 12'h333;
			{8'd126, 8'd106}: color_data = 12'h333;
			{8'd126, 8'd107}: color_data = 12'h333;
			{8'd126, 8'd108}: color_data = 12'h222;
			{8'd126, 8'd109}: color_data = 12'h222;
			{8'd126, 8'd110}: color_data = 12'h222;
			{8'd126, 8'd111}: color_data = 12'h222;
			{8'd126, 8'd112}: color_data = 12'h222;
			{8'd126, 8'd113}: color_data = 12'h222;
			{8'd126, 8'd114}: color_data = 12'h222;
			{8'd126, 8'd115}: color_data = 12'h222;
			{8'd126, 8'd116}: color_data = 12'h222;
			{8'd126, 8'd117}: color_data = 12'h222;
			{8'd126, 8'd118}: color_data = 12'h222;
			{8'd126, 8'd119}: color_data = 12'h532;
			{8'd126, 8'd120}: color_data = 12'ha23;
			{8'd126, 8'd121}: color_data = 12'hb34;
			{8'd126, 8'd122}: color_data = 12'hb56;
			{8'd126, 8'd123}: color_data = 12'hc78;
			{8'd126, 8'd124}: color_data = 12'h744;
			{8'd126, 8'd125}: color_data = 12'h432;
			{8'd126, 8'd126}: color_data = 12'h543;
			{8'd126, 8'd127}: color_data = 12'h764;
			{8'd126, 8'd128}: color_data = 12'hc96;
			{8'd126, 8'd129}: color_data = 12'h433;
			{8'd126, 8'd130}: color_data = 12'h444;
			{8'd126, 8'd131}: color_data = 12'hddd;
			{8'd126, 8'd132}: color_data = 12'hfff;
			{8'd126, 8'd133}: color_data = 12'hfff;
			{8'd126, 8'd134}: color_data = 12'hfff;
			{8'd126, 8'd135}: color_data = 12'hfff;
			{8'd126, 8'd136}: color_data = 12'hfff;
			{8'd126, 8'd137}: color_data = 12'hfff;
			{8'd126, 8'd138}: color_data = 12'hfff;
			{8'd126, 8'd139}: color_data = 12'hfff;
			{8'd126, 8'd140}: color_data = 12'hbbb;
			{8'd126, 8'd141}: color_data = 12'h777;
			{8'd127, 8'd0}: color_data = 12'hbbb;
			{8'd127, 8'd1}: color_data = 12'hbbb;
			{8'd127, 8'd2}: color_data = 12'hbbb;
			{8'd127, 8'd3}: color_data = 12'hbbb;
			{8'd127, 8'd4}: color_data = 12'haaa;
			{8'd127, 8'd5}: color_data = 12'haaa;
			{8'd127, 8'd6}: color_data = 12'haaa;
			{8'd127, 8'd7}: color_data = 12'haaa;
			{8'd127, 8'd8}: color_data = 12'haaa;
			{8'd127, 8'd9}: color_data = 12'haaa;
			{8'd127, 8'd10}: color_data = 12'haaa;
			{8'd127, 8'd11}: color_data = 12'haaa;
			{8'd127, 8'd12}: color_data = 12'haaa;
			{8'd127, 8'd13}: color_data = 12'haaa;
			{8'd127, 8'd14}: color_data = 12'haaa;
			{8'd127, 8'd15}: color_data = 12'haaa;
			{8'd127, 8'd16}: color_data = 12'haaa;
			{8'd127, 8'd17}: color_data = 12'h999;
			{8'd127, 8'd18}: color_data = 12'h999;
			{8'd127, 8'd19}: color_data = 12'h999;
			{8'd127, 8'd20}: color_data = 12'h999;
			{8'd127, 8'd21}: color_data = 12'h999;
			{8'd127, 8'd22}: color_data = 12'h999;
			{8'd127, 8'd23}: color_data = 12'h999;
			{8'd127, 8'd24}: color_data = 12'h999;
			{8'd127, 8'd25}: color_data = 12'h999;
			{8'd127, 8'd26}: color_data = 12'h999;
			{8'd127, 8'd27}: color_data = 12'h999;
			{8'd127, 8'd28}: color_data = 12'h999;
			{8'd127, 8'd29}: color_data = 12'h999;
			{8'd127, 8'd30}: color_data = 12'h888;
			{8'd127, 8'd31}: color_data = 12'h888;
			{8'd127, 8'd32}: color_data = 12'h888;
			{8'd127, 8'd33}: color_data = 12'h888;
			{8'd127, 8'd34}: color_data = 12'h888;
			{8'd127, 8'd35}: color_data = 12'h888;
			{8'd127, 8'd36}: color_data = 12'h888;
			{8'd127, 8'd37}: color_data = 12'h888;
			{8'd127, 8'd38}: color_data = 12'h888;
			{8'd127, 8'd39}: color_data = 12'h777;
			{8'd127, 8'd40}: color_data = 12'h777;
			{8'd127, 8'd41}: color_data = 12'h777;
			{8'd127, 8'd42}: color_data = 12'h777;
			{8'd127, 8'd43}: color_data = 12'h777;
			{8'd127, 8'd44}: color_data = 12'h777;
			{8'd127, 8'd45}: color_data = 12'h777;
			{8'd127, 8'd46}: color_data = 12'h777;
			{8'd127, 8'd47}: color_data = 12'h777;
			{8'd127, 8'd48}: color_data = 12'h777;
			{8'd127, 8'd49}: color_data = 12'h777;
			{8'd127, 8'd50}: color_data = 12'h777;
			{8'd127, 8'd51}: color_data = 12'h777;
			{8'd127, 8'd52}: color_data = 12'h777;
			{8'd127, 8'd53}: color_data = 12'h777;
			{8'd127, 8'd54}: color_data = 12'h777;
			{8'd127, 8'd55}: color_data = 12'h777;
			{8'd127, 8'd56}: color_data = 12'h666;
			{8'd127, 8'd57}: color_data = 12'h666;
			{8'd127, 8'd58}: color_data = 12'h666;
			{8'd127, 8'd59}: color_data = 12'h666;
			{8'd127, 8'd60}: color_data = 12'h666;
			{8'd127, 8'd61}: color_data = 12'h666;
			{8'd127, 8'd62}: color_data = 12'h666;
			{8'd127, 8'd63}: color_data = 12'h666;
			{8'd127, 8'd64}: color_data = 12'h666;
			{8'd127, 8'd65}: color_data = 12'h666;
			{8'd127, 8'd66}: color_data = 12'h666;
			{8'd127, 8'd67}: color_data = 12'h666;
			{8'd127, 8'd68}: color_data = 12'h666;
			{8'd127, 8'd69}: color_data = 12'h555;
			{8'd127, 8'd70}: color_data = 12'h555;
			{8'd127, 8'd71}: color_data = 12'h555;
			{8'd127, 8'd72}: color_data = 12'h555;
			{8'd127, 8'd73}: color_data = 12'h555;
			{8'd127, 8'd74}: color_data = 12'h555;
			{8'd127, 8'd75}: color_data = 12'h555;
			{8'd127, 8'd76}: color_data = 12'h555;
			{8'd127, 8'd77}: color_data = 12'h555;
			{8'd127, 8'd78}: color_data = 12'h555;
			{8'd127, 8'd79}: color_data = 12'h555;
			{8'd127, 8'd80}: color_data = 12'h555;
			{8'd127, 8'd81}: color_data = 12'h555;
			{8'd127, 8'd82}: color_data = 12'h444;
			{8'd127, 8'd83}: color_data = 12'h444;
			{8'd127, 8'd84}: color_data = 12'h444;
			{8'd127, 8'd85}: color_data = 12'h444;
			{8'd127, 8'd86}: color_data = 12'h444;
			{8'd127, 8'd87}: color_data = 12'h444;
			{8'd127, 8'd88}: color_data = 12'h444;
			{8'd127, 8'd89}: color_data = 12'h444;
			{8'd127, 8'd90}: color_data = 12'h444;
			{8'd127, 8'd91}: color_data = 12'h444;
			{8'd127, 8'd92}: color_data = 12'h444;
			{8'd127, 8'd93}: color_data = 12'h444;
			{8'd127, 8'd94}: color_data = 12'h444;
			{8'd127, 8'd95}: color_data = 12'h333;
			{8'd127, 8'd96}: color_data = 12'h333;
			{8'd127, 8'd97}: color_data = 12'h333;
			{8'd127, 8'd98}: color_data = 12'h333;
			{8'd127, 8'd99}: color_data = 12'h333;
			{8'd127, 8'd100}: color_data = 12'h333;
			{8'd127, 8'd101}: color_data = 12'h333;
			{8'd127, 8'd102}: color_data = 12'h333;
			{8'd127, 8'd103}: color_data = 12'h333;
			{8'd127, 8'd104}: color_data = 12'h333;
			{8'd127, 8'd105}: color_data = 12'h333;
			{8'd127, 8'd106}: color_data = 12'h333;
			{8'd127, 8'd107}: color_data = 12'h333;
			{8'd127, 8'd108}: color_data = 12'h222;
			{8'd127, 8'd109}: color_data = 12'h222;
			{8'd127, 8'd110}: color_data = 12'h222;
			{8'd127, 8'd111}: color_data = 12'h222;
			{8'd127, 8'd112}: color_data = 12'h222;
			{8'd127, 8'd113}: color_data = 12'h222;
			{8'd127, 8'd114}: color_data = 12'h222;
			{8'd127, 8'd115}: color_data = 12'h222;
			{8'd127, 8'd116}: color_data = 12'h222;
			{8'd127, 8'd117}: color_data = 12'h222;
			{8'd127, 8'd118}: color_data = 12'h222;
			{8'd127, 8'd119}: color_data = 12'h532;
			{8'd127, 8'd120}: color_data = 12'ha23;
			{8'd127, 8'd121}: color_data = 12'hb45;
			{8'd127, 8'd122}: color_data = 12'hbaa;
			{8'd127, 8'd123}: color_data = 12'ha99;
			{8'd127, 8'd124}: color_data = 12'h544;
			{8'd127, 8'd125}: color_data = 12'h432;
			{8'd127, 8'd126}: color_data = 12'h864;
			{8'd127, 8'd127}: color_data = 12'ha75;
			{8'd127, 8'd128}: color_data = 12'hc96;
			{8'd127, 8'd129}: color_data = 12'h864;
			{8'd127, 8'd130}: color_data = 12'h544;
			{8'd127, 8'd131}: color_data = 12'heee;
			{8'd127, 8'd132}: color_data = 12'hfff;
			{8'd127, 8'd133}: color_data = 12'hfff;
			{8'd127, 8'd134}: color_data = 12'hfff;
			{8'd127, 8'd135}: color_data = 12'hfff;
			{8'd127, 8'd136}: color_data = 12'hfff;
			{8'd127, 8'd137}: color_data = 12'hfff;
			{8'd127, 8'd138}: color_data = 12'hfff;
			{8'd127, 8'd139}: color_data = 12'hfff;
			{8'd127, 8'd140}: color_data = 12'haaa;
			{8'd127, 8'd141}: color_data = 12'h666;
			{8'd128, 8'd0}: color_data = 12'hbbb;
			{8'd128, 8'd1}: color_data = 12'hbbb;
			{8'd128, 8'd2}: color_data = 12'hbbb;
			{8'd128, 8'd3}: color_data = 12'hbbb;
			{8'd128, 8'd4}: color_data = 12'hbbb;
			{8'd128, 8'd5}: color_data = 12'hbbb;
			{8'd128, 8'd6}: color_data = 12'haaa;
			{8'd128, 8'd7}: color_data = 12'haaa;
			{8'd128, 8'd8}: color_data = 12'haaa;
			{8'd128, 8'd9}: color_data = 12'haaa;
			{8'd128, 8'd10}: color_data = 12'haaa;
			{8'd128, 8'd11}: color_data = 12'haaa;
			{8'd128, 8'd12}: color_data = 12'haaa;
			{8'd128, 8'd13}: color_data = 12'haaa;
			{8'd128, 8'd14}: color_data = 12'haaa;
			{8'd128, 8'd15}: color_data = 12'haaa;
			{8'd128, 8'd16}: color_data = 12'haaa;
			{8'd128, 8'd17}: color_data = 12'h999;
			{8'd128, 8'd18}: color_data = 12'h999;
			{8'd128, 8'd19}: color_data = 12'h999;
			{8'd128, 8'd20}: color_data = 12'h999;
			{8'd128, 8'd21}: color_data = 12'h999;
			{8'd128, 8'd22}: color_data = 12'h999;
			{8'd128, 8'd23}: color_data = 12'h999;
			{8'd128, 8'd24}: color_data = 12'h999;
			{8'd128, 8'd25}: color_data = 12'h999;
			{8'd128, 8'd26}: color_data = 12'h999;
			{8'd128, 8'd27}: color_data = 12'h999;
			{8'd128, 8'd28}: color_data = 12'h999;
			{8'd128, 8'd29}: color_data = 12'h999;
			{8'd128, 8'd30}: color_data = 12'h888;
			{8'd128, 8'd31}: color_data = 12'h888;
			{8'd128, 8'd32}: color_data = 12'h888;
			{8'd128, 8'd33}: color_data = 12'h888;
			{8'd128, 8'd34}: color_data = 12'h888;
			{8'd128, 8'd35}: color_data = 12'h888;
			{8'd128, 8'd36}: color_data = 12'h888;
			{8'd128, 8'd37}: color_data = 12'h888;
			{8'd128, 8'd38}: color_data = 12'h777;
			{8'd128, 8'd39}: color_data = 12'h566;
			{8'd128, 8'd40}: color_data = 12'h456;
			{8'd128, 8'd41}: color_data = 12'h678;
			{8'd128, 8'd42}: color_data = 12'h678;
			{8'd128, 8'd43}: color_data = 12'h677;
			{8'd128, 8'd44}: color_data = 12'h677;
			{8'd128, 8'd45}: color_data = 12'h577;
			{8'd128, 8'd46}: color_data = 12'h678;
			{8'd128, 8'd47}: color_data = 12'h777;
			{8'd128, 8'd48}: color_data = 12'h777;
			{8'd128, 8'd49}: color_data = 12'h777;
			{8'd128, 8'd50}: color_data = 12'h777;
			{8'd128, 8'd51}: color_data = 12'h777;
			{8'd128, 8'd52}: color_data = 12'h777;
			{8'd128, 8'd53}: color_data = 12'h777;
			{8'd128, 8'd54}: color_data = 12'h777;
			{8'd128, 8'd55}: color_data = 12'h777;
			{8'd128, 8'd56}: color_data = 12'h666;
			{8'd128, 8'd57}: color_data = 12'h666;
			{8'd128, 8'd58}: color_data = 12'h666;
			{8'd128, 8'd59}: color_data = 12'h666;
			{8'd128, 8'd60}: color_data = 12'h666;
			{8'd128, 8'd61}: color_data = 12'h666;
			{8'd128, 8'd62}: color_data = 12'h666;
			{8'd128, 8'd63}: color_data = 12'h666;
			{8'd128, 8'd64}: color_data = 12'h666;
			{8'd128, 8'd65}: color_data = 12'h666;
			{8'd128, 8'd66}: color_data = 12'h666;
			{8'd128, 8'd67}: color_data = 12'h666;
			{8'd128, 8'd68}: color_data = 12'h666;
			{8'd128, 8'd69}: color_data = 12'h555;
			{8'd128, 8'd70}: color_data = 12'h555;
			{8'd128, 8'd71}: color_data = 12'h555;
			{8'd128, 8'd72}: color_data = 12'h555;
			{8'd128, 8'd73}: color_data = 12'h555;
			{8'd128, 8'd74}: color_data = 12'h555;
			{8'd128, 8'd75}: color_data = 12'h555;
			{8'd128, 8'd76}: color_data = 12'h555;
			{8'd128, 8'd77}: color_data = 12'h555;
			{8'd128, 8'd78}: color_data = 12'h555;
			{8'd128, 8'd79}: color_data = 12'h555;
			{8'd128, 8'd80}: color_data = 12'h555;
			{8'd128, 8'd81}: color_data = 12'h555;
			{8'd128, 8'd82}: color_data = 12'h444;
			{8'd128, 8'd83}: color_data = 12'h444;
			{8'd128, 8'd84}: color_data = 12'h444;
			{8'd128, 8'd85}: color_data = 12'h444;
			{8'd128, 8'd86}: color_data = 12'h444;
			{8'd128, 8'd87}: color_data = 12'h444;
			{8'd128, 8'd88}: color_data = 12'h444;
			{8'd128, 8'd89}: color_data = 12'h444;
			{8'd128, 8'd90}: color_data = 12'h444;
			{8'd128, 8'd91}: color_data = 12'h444;
			{8'd128, 8'd92}: color_data = 12'h444;
			{8'd128, 8'd93}: color_data = 12'h444;
			{8'd128, 8'd94}: color_data = 12'h444;
			{8'd128, 8'd95}: color_data = 12'h333;
			{8'd128, 8'd96}: color_data = 12'h333;
			{8'd128, 8'd97}: color_data = 12'h333;
			{8'd128, 8'd98}: color_data = 12'h333;
			{8'd128, 8'd99}: color_data = 12'h333;
			{8'd128, 8'd100}: color_data = 12'h333;
			{8'd128, 8'd101}: color_data = 12'h333;
			{8'd128, 8'd102}: color_data = 12'h333;
			{8'd128, 8'd103}: color_data = 12'h333;
			{8'd128, 8'd104}: color_data = 12'h333;
			{8'd128, 8'd105}: color_data = 12'h333;
			{8'd128, 8'd106}: color_data = 12'h333;
			{8'd128, 8'd107}: color_data = 12'h333;
			{8'd128, 8'd108}: color_data = 12'h222;
			{8'd128, 8'd109}: color_data = 12'h222;
			{8'd128, 8'd110}: color_data = 12'h222;
			{8'd128, 8'd111}: color_data = 12'h222;
			{8'd128, 8'd112}: color_data = 12'h222;
			{8'd128, 8'd113}: color_data = 12'h222;
			{8'd128, 8'd114}: color_data = 12'h222;
			{8'd128, 8'd115}: color_data = 12'h222;
			{8'd128, 8'd116}: color_data = 12'h222;
			{8'd128, 8'd117}: color_data = 12'h222;
			{8'd128, 8'd118}: color_data = 12'h222;
			{8'd128, 8'd119}: color_data = 12'h422;
			{8'd128, 8'd120}: color_data = 12'h822;
			{8'd128, 8'd121}: color_data = 12'hb55;
			{8'd128, 8'd122}: color_data = 12'hbbb;
			{8'd128, 8'd123}: color_data = 12'h844;
			{8'd128, 8'd124}: color_data = 12'h422;
			{8'd128, 8'd125}: color_data = 12'h432;
			{8'd128, 8'd126}: color_data = 12'h864;
			{8'd128, 8'd127}: color_data = 12'hb85;
			{8'd128, 8'd128}: color_data = 12'hc96;
			{8'd128, 8'd129}: color_data = 12'hb85;
			{8'd128, 8'd130}: color_data = 12'h655;
			{8'd128, 8'd131}: color_data = 12'heff;
			{8'd128, 8'd132}: color_data = 12'hfff;
			{8'd128, 8'd133}: color_data = 12'hfff;
			{8'd128, 8'd134}: color_data = 12'hfff;
			{8'd128, 8'd135}: color_data = 12'hfff;
			{8'd128, 8'd136}: color_data = 12'hfff;
			{8'd128, 8'd137}: color_data = 12'hfff;
			{8'd128, 8'd138}: color_data = 12'hfff;
			{8'd128, 8'd139}: color_data = 12'hfff;
			{8'd128, 8'd140}: color_data = 12'haaa;
			{8'd128, 8'd141}: color_data = 12'h555;
			{8'd129, 8'd0}: color_data = 12'hbbb;
			{8'd129, 8'd1}: color_data = 12'hbbb;
			{8'd129, 8'd2}: color_data = 12'hbbb;
			{8'd129, 8'd3}: color_data = 12'hbbb;
			{8'd129, 8'd4}: color_data = 12'haaa;
			{8'd129, 8'd5}: color_data = 12'haaa;
			{8'd129, 8'd6}: color_data = 12'haaa;
			{8'd129, 8'd7}: color_data = 12'haaa;
			{8'd129, 8'd8}: color_data = 12'hbbb;
			{8'd129, 8'd9}: color_data = 12'haaa;
			{8'd129, 8'd10}: color_data = 12'haaa;
			{8'd129, 8'd11}: color_data = 12'haaa;
			{8'd129, 8'd12}: color_data = 12'haaa;
			{8'd129, 8'd13}: color_data = 12'haaa;
			{8'd129, 8'd14}: color_data = 12'haaa;
			{8'd129, 8'd15}: color_data = 12'haaa;
			{8'd129, 8'd16}: color_data = 12'haaa;
			{8'd129, 8'd17}: color_data = 12'h999;
			{8'd129, 8'd18}: color_data = 12'h999;
			{8'd129, 8'd19}: color_data = 12'h999;
			{8'd129, 8'd20}: color_data = 12'h999;
			{8'd129, 8'd21}: color_data = 12'h999;
			{8'd129, 8'd22}: color_data = 12'h999;
			{8'd129, 8'd23}: color_data = 12'h999;
			{8'd129, 8'd24}: color_data = 12'h999;
			{8'd129, 8'd25}: color_data = 12'h999;
			{8'd129, 8'd26}: color_data = 12'h999;
			{8'd129, 8'd27}: color_data = 12'h999;
			{8'd129, 8'd28}: color_data = 12'h999;
			{8'd129, 8'd29}: color_data = 12'h999;
			{8'd129, 8'd30}: color_data = 12'h888;
			{8'd129, 8'd31}: color_data = 12'h888;
			{8'd129, 8'd32}: color_data = 12'h888;
			{8'd129, 8'd33}: color_data = 12'h888;
			{8'd129, 8'd34}: color_data = 12'h888;
			{8'd129, 8'd35}: color_data = 12'h888;
			{8'd129, 8'd36}: color_data = 12'h888;
			{8'd129, 8'd37}: color_data = 12'h888;
			{8'd129, 8'd38}: color_data = 12'h455;
			{8'd129, 8'd39}: color_data = 12'hb20;
			{8'd129, 8'd40}: color_data = 12'hb30;
			{8'd129, 8'd41}: color_data = 12'ha40;
			{8'd129, 8'd42}: color_data = 12'ha40;
			{8'd129, 8'd43}: color_data = 12'ha40;
			{8'd129, 8'd44}: color_data = 12'ha40;
			{8'd129, 8'd45}: color_data = 12'hb50;
			{8'd129, 8'd46}: color_data = 12'ha50;
			{8'd129, 8'd48}: color_data = 12'h677;
			{8'd129, 8'd49}: color_data = 12'h777;
			{8'd129, 8'd50}: color_data = 12'h777;
			{8'd129, 8'd51}: color_data = 12'h777;
			{8'd129, 8'd52}: color_data = 12'h777;
			{8'd129, 8'd53}: color_data = 12'h777;
			{8'd129, 8'd54}: color_data = 12'h777;
			{8'd129, 8'd55}: color_data = 12'h777;
			{8'd129, 8'd56}: color_data = 12'h666;
			{8'd129, 8'd57}: color_data = 12'h666;
			{8'd129, 8'd58}: color_data = 12'h666;
			{8'd129, 8'd59}: color_data = 12'h666;
			{8'd129, 8'd60}: color_data = 12'h666;
			{8'd129, 8'd61}: color_data = 12'h666;
			{8'd129, 8'd62}: color_data = 12'h666;
			{8'd129, 8'd63}: color_data = 12'h666;
			{8'd129, 8'd64}: color_data = 12'h666;
			{8'd129, 8'd65}: color_data = 12'h666;
			{8'd129, 8'd66}: color_data = 12'h666;
			{8'd129, 8'd67}: color_data = 12'h666;
			{8'd129, 8'd68}: color_data = 12'h666;
			{8'd129, 8'd69}: color_data = 12'h555;
			{8'd129, 8'd70}: color_data = 12'h555;
			{8'd129, 8'd71}: color_data = 12'h555;
			{8'd129, 8'd72}: color_data = 12'h555;
			{8'd129, 8'd73}: color_data = 12'h555;
			{8'd129, 8'd74}: color_data = 12'h555;
			{8'd129, 8'd75}: color_data = 12'h555;
			{8'd129, 8'd76}: color_data = 12'h555;
			{8'd129, 8'd77}: color_data = 12'h555;
			{8'd129, 8'd78}: color_data = 12'h555;
			{8'd129, 8'd79}: color_data = 12'h555;
			{8'd129, 8'd80}: color_data = 12'h555;
			{8'd129, 8'd81}: color_data = 12'h555;
			{8'd129, 8'd82}: color_data = 12'h444;
			{8'd129, 8'd83}: color_data = 12'h444;
			{8'd129, 8'd84}: color_data = 12'h444;
			{8'd129, 8'd85}: color_data = 12'h444;
			{8'd129, 8'd86}: color_data = 12'h444;
			{8'd129, 8'd87}: color_data = 12'h444;
			{8'd129, 8'd88}: color_data = 12'h444;
			{8'd129, 8'd89}: color_data = 12'h444;
			{8'd129, 8'd90}: color_data = 12'h444;
			{8'd129, 8'd91}: color_data = 12'h444;
			{8'd129, 8'd92}: color_data = 12'h444;
			{8'd129, 8'd93}: color_data = 12'h444;
			{8'd129, 8'd94}: color_data = 12'h444;
			{8'd129, 8'd95}: color_data = 12'h333;
			{8'd129, 8'd96}: color_data = 12'h333;
			{8'd129, 8'd97}: color_data = 12'h333;
			{8'd129, 8'd98}: color_data = 12'h333;
			{8'd129, 8'd99}: color_data = 12'h333;
			{8'd129, 8'd100}: color_data = 12'h333;
			{8'd129, 8'd101}: color_data = 12'h333;
			{8'd129, 8'd102}: color_data = 12'h333;
			{8'd129, 8'd103}: color_data = 12'h333;
			{8'd129, 8'd104}: color_data = 12'h333;
			{8'd129, 8'd105}: color_data = 12'h333;
			{8'd129, 8'd106}: color_data = 12'h333;
			{8'd129, 8'd107}: color_data = 12'h333;
			{8'd129, 8'd108}: color_data = 12'h222;
			{8'd129, 8'd109}: color_data = 12'h222;
			{8'd129, 8'd110}: color_data = 12'h222;
			{8'd129, 8'd111}: color_data = 12'h222;
			{8'd129, 8'd112}: color_data = 12'h222;
			{8'd129, 8'd113}: color_data = 12'h222;
			{8'd129, 8'd114}: color_data = 12'h222;
			{8'd129, 8'd115}: color_data = 12'h222;
			{8'd129, 8'd116}: color_data = 12'h222;
			{8'd129, 8'd117}: color_data = 12'h222;
			{8'd129, 8'd118}: color_data = 12'h222;
			{8'd129, 8'd119}: color_data = 12'h222;
			{8'd129, 8'd120}: color_data = 12'h622;
			{8'd129, 8'd121}: color_data = 12'h933;
			{8'd129, 8'd122}: color_data = 12'hb77;
			{8'd129, 8'd123}: color_data = 12'ha66;
			{8'd129, 8'd124}: color_data = 12'h544;
			{8'd129, 8'd125}: color_data = 12'h322;
			{8'd129, 8'd126}: color_data = 12'h643;
			{8'd129, 8'd127}: color_data = 12'hb85;
			{8'd129, 8'd128}: color_data = 12'hc96;
			{8'd129, 8'd129}: color_data = 12'hb85;
			{8'd129, 8'd130}: color_data = 12'h765;
			{8'd129, 8'd131}: color_data = 12'hfff;
			{8'd129, 8'd132}: color_data = 12'hfff;
			{8'd129, 8'd133}: color_data = 12'hfff;
			{8'd129, 8'd134}: color_data = 12'hfff;
			{8'd129, 8'd135}: color_data = 12'hfff;
			{8'd129, 8'd136}: color_data = 12'hfff;
			{8'd129, 8'd137}: color_data = 12'hfff;
			{8'd129, 8'd138}: color_data = 12'hfff;
			{8'd129, 8'd139}: color_data = 12'heee;
			{8'd129, 8'd140}: color_data = 12'haaa;
			{8'd129, 8'd141}: color_data = 12'h333;
			{8'd130, 8'd2}: color_data = 12'hfff;
			{8'd130, 8'd3}: color_data = 12'hbbb;
			{8'd130, 8'd4}: color_data = 12'haaa;
			{8'd130, 8'd5}: color_data = 12'hbbb;
			{8'd130, 8'd6}: color_data = 12'haaa;
			{8'd130, 8'd7}: color_data = 12'haaa;
			{8'd130, 8'd8}: color_data = 12'haaa;
			{8'd130, 8'd9}: color_data = 12'haaa;
			{8'd130, 8'd10}: color_data = 12'haaa;
			{8'd130, 8'd11}: color_data = 12'haaa;
			{8'd130, 8'd12}: color_data = 12'haaa;
			{8'd130, 8'd13}: color_data = 12'haaa;
			{8'd130, 8'd14}: color_data = 12'haaa;
			{8'd130, 8'd15}: color_data = 12'haaa;
			{8'd130, 8'd16}: color_data = 12'haaa;
			{8'd130, 8'd17}: color_data = 12'haaa;
			{8'd130, 8'd18}: color_data = 12'h999;
			{8'd130, 8'd19}: color_data = 12'h999;
			{8'd130, 8'd20}: color_data = 12'h999;
			{8'd130, 8'd21}: color_data = 12'h999;
			{8'd130, 8'd22}: color_data = 12'h999;
			{8'd130, 8'd23}: color_data = 12'h999;
			{8'd130, 8'd24}: color_data = 12'h999;
			{8'd130, 8'd25}: color_data = 12'h999;
			{8'd130, 8'd26}: color_data = 12'h999;
			{8'd130, 8'd27}: color_data = 12'h999;
			{8'd130, 8'd28}: color_data = 12'h999;
			{8'd130, 8'd29}: color_data = 12'h999;
			{8'd130, 8'd30}: color_data = 12'h888;
			{8'd130, 8'd31}: color_data = 12'h888;
			{8'd130, 8'd32}: color_data = 12'h888;
			{8'd130, 8'd33}: color_data = 12'h888;
			{8'd130, 8'd34}: color_data = 12'h888;
			{8'd130, 8'd35}: color_data = 12'h888;
			{8'd130, 8'd36}: color_data = 12'h888;
			{8'd130, 8'd37}: color_data = 12'h7ff;
			{8'd130, 8'd38}: color_data = 12'ha20;
			{8'd130, 8'd39}: color_data = 12'hc41;
			{8'd130, 8'd40}: color_data = 12'hc41;
			{8'd130, 8'd41}: color_data = 12'hc51;
			{8'd130, 8'd42}: color_data = 12'hc51;
			{8'd130, 8'd43}: color_data = 12'hc51;
			{8'd130, 8'd44}: color_data = 12'hc61;
			{8'd130, 8'd45}: color_data = 12'hc61;
			{8'd130, 8'd46}: color_data = 12'hc61;
			{8'd130, 8'd47}: color_data = 12'hc60;
			{8'd130, 8'd48}: color_data = 12'hb60;
			{8'd130, 8'd49}: color_data = 12'h667;
			{8'd130, 8'd50}: color_data = 12'h677;
			{8'd130, 8'd51}: color_data = 12'h777;
			{8'd130, 8'd52}: color_data = 12'h777;
			{8'd130, 8'd53}: color_data = 12'h777;
			{8'd130, 8'd54}: color_data = 12'h777;
			{8'd130, 8'd55}: color_data = 12'h777;
			{8'd130, 8'd56}: color_data = 12'h666;
			{8'd130, 8'd57}: color_data = 12'h666;
			{8'd130, 8'd58}: color_data = 12'h666;
			{8'd130, 8'd59}: color_data = 12'h666;
			{8'd130, 8'd60}: color_data = 12'h666;
			{8'd130, 8'd61}: color_data = 12'h666;
			{8'd130, 8'd62}: color_data = 12'h666;
			{8'd130, 8'd63}: color_data = 12'h666;
			{8'd130, 8'd64}: color_data = 12'h666;
			{8'd130, 8'd65}: color_data = 12'h666;
			{8'd130, 8'd66}: color_data = 12'h666;
			{8'd130, 8'd67}: color_data = 12'h666;
			{8'd130, 8'd68}: color_data = 12'h666;
			{8'd130, 8'd69}: color_data = 12'h555;
			{8'd130, 8'd70}: color_data = 12'h555;
			{8'd130, 8'd71}: color_data = 12'h555;
			{8'd130, 8'd72}: color_data = 12'h555;
			{8'd130, 8'd73}: color_data = 12'h555;
			{8'd130, 8'd74}: color_data = 12'h555;
			{8'd130, 8'd75}: color_data = 12'h555;
			{8'd130, 8'd76}: color_data = 12'h555;
			{8'd130, 8'd77}: color_data = 12'h555;
			{8'd130, 8'd78}: color_data = 12'h555;
			{8'd130, 8'd79}: color_data = 12'h555;
			{8'd130, 8'd80}: color_data = 12'h555;
			{8'd130, 8'd81}: color_data = 12'h555;
			{8'd130, 8'd82}: color_data = 12'h444;
			{8'd130, 8'd83}: color_data = 12'h444;
			{8'd130, 8'd84}: color_data = 12'h444;
			{8'd130, 8'd85}: color_data = 12'h444;
			{8'd130, 8'd86}: color_data = 12'h444;
			{8'd130, 8'd87}: color_data = 12'h444;
			{8'd130, 8'd88}: color_data = 12'h444;
			{8'd130, 8'd89}: color_data = 12'h444;
			{8'd130, 8'd90}: color_data = 12'h444;
			{8'd130, 8'd91}: color_data = 12'h444;
			{8'd130, 8'd92}: color_data = 12'h444;
			{8'd130, 8'd93}: color_data = 12'h444;
			{8'd130, 8'd94}: color_data = 12'h444;
			{8'd130, 8'd95}: color_data = 12'h333;
			{8'd130, 8'd96}: color_data = 12'h333;
			{8'd130, 8'd97}: color_data = 12'h333;
			{8'd130, 8'd98}: color_data = 12'h333;
			{8'd130, 8'd99}: color_data = 12'h333;
			{8'd130, 8'd100}: color_data = 12'h333;
			{8'd130, 8'd101}: color_data = 12'h333;
			{8'd130, 8'd102}: color_data = 12'h333;
			{8'd130, 8'd103}: color_data = 12'h333;
			{8'd130, 8'd104}: color_data = 12'h333;
			{8'd130, 8'd105}: color_data = 12'h333;
			{8'd130, 8'd106}: color_data = 12'h333;
			{8'd130, 8'd107}: color_data = 12'h333;
			{8'd130, 8'd108}: color_data = 12'h222;
			{8'd130, 8'd109}: color_data = 12'h222;
			{8'd130, 8'd110}: color_data = 12'h222;
			{8'd130, 8'd111}: color_data = 12'h222;
			{8'd130, 8'd112}: color_data = 12'h222;
			{8'd130, 8'd113}: color_data = 12'h222;
			{8'd130, 8'd114}: color_data = 12'h222;
			{8'd130, 8'd115}: color_data = 12'h222;
			{8'd130, 8'd116}: color_data = 12'h222;
			{8'd130, 8'd117}: color_data = 12'h222;
			{8'd130, 8'd118}: color_data = 12'h222;
			{8'd130, 8'd119}: color_data = 12'h222;
			{8'd130, 8'd120}: color_data = 12'h322;
			{8'd130, 8'd121}: color_data = 12'h522;
			{8'd130, 8'd122}: color_data = 12'h722;
			{8'd130, 8'd123}: color_data = 12'h722;
			{8'd130, 8'd124}: color_data = 12'h322;
			{8'd130, 8'd125}: color_data = 12'h322;
			{8'd130, 8'd126}: color_data = 12'h864;
			{8'd130, 8'd127}: color_data = 12'hc96;
			{8'd130, 8'd128}: color_data = 12'hc96;
			{8'd130, 8'd129}: color_data = 12'ha85;
			{8'd130, 8'd130}: color_data = 12'h765;
			{8'd130, 8'd131}: color_data = 12'hfff;
			{8'd130, 8'd132}: color_data = 12'hfff;
			{8'd130, 8'd133}: color_data = 12'hfff;
			{8'd130, 8'd134}: color_data = 12'hfff;
			{8'd130, 8'd135}: color_data = 12'hfff;
			{8'd130, 8'd136}: color_data = 12'hfff;
			{8'd130, 8'd137}: color_data = 12'hfff;
			{8'd130, 8'd138}: color_data = 12'hfff;
			{8'd130, 8'd139}: color_data = 12'heee;
			{8'd130, 8'd140}: color_data = 12'h999;
			{8'd130, 8'd141}: color_data = 12'h555;
			{8'd131, 8'd7}: color_data = 12'h777;
			{8'd131, 8'd8}: color_data = 12'hbbb;
			{8'd131, 8'd9}: color_data = 12'h999;
			{8'd131, 8'd10}: color_data = 12'haaa;
			{8'd131, 8'd11}: color_data = 12'haaa;
			{8'd131, 8'd12}: color_data = 12'haaa;
			{8'd131, 8'd13}: color_data = 12'haaa;
			{8'd131, 8'd14}: color_data = 12'haaa;
			{8'd131, 8'd15}: color_data = 12'haaa;
			{8'd131, 8'd16}: color_data = 12'haaa;
			{8'd131, 8'd17}: color_data = 12'haaa;
			{8'd131, 8'd18}: color_data = 12'haaa;
			{8'd131, 8'd19}: color_data = 12'haaa;
			{8'd131, 8'd20}: color_data = 12'ha99;
			{8'd131, 8'd21}: color_data = 12'h999;
			{8'd131, 8'd22}: color_data = 12'h999;
			{8'd131, 8'd23}: color_data = 12'h999;
			{8'd131, 8'd24}: color_data = 12'h999;
			{8'd131, 8'd25}: color_data = 12'h999;
			{8'd131, 8'd26}: color_data = 12'h999;
			{8'd131, 8'd27}: color_data = 12'h999;
			{8'd131, 8'd28}: color_data = 12'h999;
			{8'd131, 8'd29}: color_data = 12'h999;
			{8'd131, 8'd30}: color_data = 12'h888;
			{8'd131, 8'd31}: color_data = 12'h888;
			{8'd131, 8'd32}: color_data = 12'h888;
			{8'd131, 8'd33}: color_data = 12'h888;
			{8'd131, 8'd34}: color_data = 12'h888;
			{8'd131, 8'd35}: color_data = 12'h888;
			{8'd131, 8'd36}: color_data = 12'h788;
			{8'd131, 8'd37}: color_data = 12'ha20;
			{8'd131, 8'd38}: color_data = 12'hc41;
			{8'd131, 8'd39}: color_data = 12'hd41;
			{8'd131, 8'd40}: color_data = 12'he51;
			{8'd131, 8'd41}: color_data = 12'he61;
			{8'd131, 8'd42}: color_data = 12'he61;
			{8'd131, 8'd43}: color_data = 12'he61;
			{8'd131, 8'd44}: color_data = 12'he71;
			{8'd131, 8'd45}: color_data = 12'he71;
			{8'd131, 8'd46}: color_data = 12'he71;
			{8'd131, 8'd47}: color_data = 12'hd70;
			{8'd131, 8'd48}: color_data = 12'hc70;
			{8'd131, 8'd49}: color_data = 12'ha50;
			{8'd131, 8'd50}: color_data = 12'h578;
			{8'd131, 8'd51}: color_data = 12'h777;
			{8'd131, 8'd52}: color_data = 12'h777;
			{8'd131, 8'd53}: color_data = 12'h777;
			{8'd131, 8'd54}: color_data = 12'h777;
			{8'd131, 8'd55}: color_data = 12'h777;
			{8'd131, 8'd56}: color_data = 12'h666;
			{8'd131, 8'd57}: color_data = 12'h666;
			{8'd131, 8'd58}: color_data = 12'h666;
			{8'd131, 8'd59}: color_data = 12'h666;
			{8'd131, 8'd60}: color_data = 12'h666;
			{8'd131, 8'd61}: color_data = 12'h666;
			{8'd131, 8'd62}: color_data = 12'h666;
			{8'd131, 8'd63}: color_data = 12'h666;
			{8'd131, 8'd64}: color_data = 12'h666;
			{8'd131, 8'd65}: color_data = 12'h666;
			{8'd131, 8'd66}: color_data = 12'h666;
			{8'd131, 8'd67}: color_data = 12'h666;
			{8'd131, 8'd68}: color_data = 12'h666;
			{8'd131, 8'd69}: color_data = 12'h555;
			{8'd131, 8'd70}: color_data = 12'h555;
			{8'd131, 8'd71}: color_data = 12'h555;
			{8'd131, 8'd72}: color_data = 12'h555;
			{8'd131, 8'd73}: color_data = 12'h555;
			{8'd131, 8'd74}: color_data = 12'h555;
			{8'd131, 8'd75}: color_data = 12'h555;
			{8'd131, 8'd76}: color_data = 12'h555;
			{8'd131, 8'd77}: color_data = 12'h555;
			{8'd131, 8'd78}: color_data = 12'h555;
			{8'd131, 8'd79}: color_data = 12'h555;
			{8'd131, 8'd80}: color_data = 12'h555;
			{8'd131, 8'd81}: color_data = 12'h555;
			{8'd131, 8'd82}: color_data = 12'h444;
			{8'd131, 8'd83}: color_data = 12'h444;
			{8'd131, 8'd84}: color_data = 12'h444;
			{8'd131, 8'd85}: color_data = 12'h444;
			{8'd131, 8'd86}: color_data = 12'h444;
			{8'd131, 8'd87}: color_data = 12'h444;
			{8'd131, 8'd88}: color_data = 12'h444;
			{8'd131, 8'd89}: color_data = 12'h444;
			{8'd131, 8'd90}: color_data = 12'h444;
			{8'd131, 8'd91}: color_data = 12'h444;
			{8'd131, 8'd92}: color_data = 12'h444;
			{8'd131, 8'd93}: color_data = 12'h444;
			{8'd131, 8'd94}: color_data = 12'h444;
			{8'd131, 8'd95}: color_data = 12'h333;
			{8'd131, 8'd96}: color_data = 12'h333;
			{8'd131, 8'd97}: color_data = 12'h333;
			{8'd131, 8'd98}: color_data = 12'h333;
			{8'd131, 8'd99}: color_data = 12'h333;
			{8'd131, 8'd100}: color_data = 12'h333;
			{8'd131, 8'd101}: color_data = 12'h333;
			{8'd131, 8'd102}: color_data = 12'h333;
			{8'd131, 8'd103}: color_data = 12'h333;
			{8'd131, 8'd104}: color_data = 12'h333;
			{8'd131, 8'd105}: color_data = 12'h333;
			{8'd131, 8'd106}: color_data = 12'h333;
			{8'd131, 8'd107}: color_data = 12'h333;
			{8'd131, 8'd108}: color_data = 12'h222;
			{8'd131, 8'd109}: color_data = 12'h222;
			{8'd131, 8'd110}: color_data = 12'h222;
			{8'd131, 8'd111}: color_data = 12'h222;
			{8'd131, 8'd112}: color_data = 12'h222;
			{8'd131, 8'd113}: color_data = 12'h222;
			{8'd131, 8'd114}: color_data = 12'h222;
			{8'd131, 8'd115}: color_data = 12'h222;
			{8'd131, 8'd116}: color_data = 12'h222;
			{8'd131, 8'd117}: color_data = 12'h222;
			{8'd131, 8'd118}: color_data = 12'h222;
			{8'd131, 8'd119}: color_data = 12'h222;
			{8'd131, 8'd120}: color_data = 12'h122;
			{8'd131, 8'd121}: color_data = 12'h222;
			{8'd131, 8'd122}: color_data = 12'h321;
			{8'd131, 8'd123}: color_data = 12'h655;
			{8'd131, 8'd124}: color_data = 12'h877;
			{8'd131, 8'd125}: color_data = 12'h222;
			{8'd131, 8'd126}: color_data = 12'h642;
			{8'd131, 8'd127}: color_data = 12'ha75;
			{8'd131, 8'd128}: color_data = 12'hb85;
			{8'd131, 8'd129}: color_data = 12'h742;
			{8'd131, 8'd130}: color_data = 12'h554;
			{8'd131, 8'd131}: color_data = 12'hfff;
			{8'd131, 8'd132}: color_data = 12'hfff;
			{8'd131, 8'd133}: color_data = 12'hfff;
			{8'd131, 8'd134}: color_data = 12'hfff;
			{8'd131, 8'd135}: color_data = 12'hfff;
			{8'd131, 8'd136}: color_data = 12'hfff;
			{8'd131, 8'd137}: color_data = 12'hfff;
			{8'd131, 8'd138}: color_data = 12'hfff;
			{8'd131, 8'd139}: color_data = 12'hddd;
			{8'd131, 8'd140}: color_data = 12'h999;
			{8'd132, 8'd13}: color_data = 12'h999;
			{8'd132, 8'd14}: color_data = 12'haaa;
			{8'd132, 8'd15}: color_data = 12'haaa;
			{8'd132, 8'd16}: color_data = 12'haaa;
			{8'd132, 8'd17}: color_data = 12'h999;
			{8'd132, 8'd18}: color_data = 12'h999;
			{8'd132, 8'd19}: color_data = 12'h999;
			{8'd132, 8'd20}: color_data = 12'h999;
			{8'd132, 8'd21}: color_data = 12'h999;
			{8'd132, 8'd22}: color_data = 12'h999;
			{8'd132, 8'd23}: color_data = 12'h999;
			{8'd132, 8'd24}: color_data = 12'h999;
			{8'd132, 8'd25}: color_data = 12'h999;
			{8'd132, 8'd26}: color_data = 12'h999;
			{8'd132, 8'd27}: color_data = 12'h999;
			{8'd132, 8'd28}: color_data = 12'h999;
			{8'd132, 8'd29}: color_data = 12'h999;
			{8'd132, 8'd30}: color_data = 12'h888;
			{8'd132, 8'd31}: color_data = 12'h888;
			{8'd132, 8'd32}: color_data = 12'h888;
			{8'd132, 8'd33}: color_data = 12'h888;
			{8'd132, 8'd34}: color_data = 12'h777;
			{8'd132, 8'd35}: color_data = 12'h69a;
			{8'd132, 8'd36}: color_data = 12'hc20;
			{8'd132, 8'd37}: color_data = 12'hd31;
			{8'd132, 8'd38}: color_data = 12'he41;
			{8'd132, 8'd39}: color_data = 12'he51;
			{8'd132, 8'd40}: color_data = 12'he51;
			{8'd132, 8'd41}: color_data = 12'he51;
			{8'd132, 8'd42}: color_data = 12'he61;
			{8'd132, 8'd43}: color_data = 12'he61;
			{8'd132, 8'd44}: color_data = 12'he71;
			{8'd132, 8'd45}: color_data = 12'he71;
			{8'd132, 8'd46}: color_data = 12'he71;
			{8'd132, 8'd47}: color_data = 12'he80;
			{8'd132, 8'd48}: color_data = 12'he80;
			{8'd132, 8'd49}: color_data = 12'hb70;
			{8'd132, 8'd50}: color_data = 12'ha60;
			{8'd132, 8'd51}: color_data = 12'h568;
			{8'd132, 8'd52}: color_data = 12'h666;
			{8'd132, 8'd53}: color_data = 12'h666;
			{8'd132, 8'd54}: color_data = 12'h777;
			{8'd132, 8'd55}: color_data = 12'h777;
			{8'd132, 8'd56}: color_data = 12'h666;
			{8'd132, 8'd57}: color_data = 12'h666;
			{8'd132, 8'd58}: color_data = 12'h666;
			{8'd132, 8'd59}: color_data = 12'h666;
			{8'd132, 8'd60}: color_data = 12'h666;
			{8'd132, 8'd61}: color_data = 12'h666;
			{8'd132, 8'd62}: color_data = 12'h666;
			{8'd132, 8'd63}: color_data = 12'h666;
			{8'd132, 8'd64}: color_data = 12'h666;
			{8'd132, 8'd65}: color_data = 12'h666;
			{8'd132, 8'd66}: color_data = 12'h666;
			{8'd132, 8'd67}: color_data = 12'h666;
			{8'd132, 8'd68}: color_data = 12'h666;
			{8'd132, 8'd69}: color_data = 12'h555;
			{8'd132, 8'd70}: color_data = 12'h555;
			{8'd132, 8'd71}: color_data = 12'h555;
			{8'd132, 8'd72}: color_data = 12'h555;
			{8'd132, 8'd73}: color_data = 12'h555;
			{8'd132, 8'd74}: color_data = 12'h555;
			{8'd132, 8'd75}: color_data = 12'h555;
			{8'd132, 8'd76}: color_data = 12'h555;
			{8'd132, 8'd77}: color_data = 12'h555;
			{8'd132, 8'd78}: color_data = 12'h555;
			{8'd132, 8'd79}: color_data = 12'h555;
			{8'd132, 8'd80}: color_data = 12'h555;
			{8'd132, 8'd81}: color_data = 12'h555;
			{8'd132, 8'd82}: color_data = 12'h444;
			{8'd132, 8'd83}: color_data = 12'h444;
			{8'd132, 8'd84}: color_data = 12'h444;
			{8'd132, 8'd85}: color_data = 12'h444;
			{8'd132, 8'd86}: color_data = 12'h444;
			{8'd132, 8'd87}: color_data = 12'h444;
			{8'd132, 8'd88}: color_data = 12'h444;
			{8'd132, 8'd89}: color_data = 12'h444;
			{8'd132, 8'd90}: color_data = 12'h444;
			{8'd132, 8'd91}: color_data = 12'h444;
			{8'd132, 8'd92}: color_data = 12'h444;
			{8'd132, 8'd93}: color_data = 12'h444;
			{8'd132, 8'd94}: color_data = 12'h444;
			{8'd132, 8'd95}: color_data = 12'h333;
			{8'd132, 8'd96}: color_data = 12'h333;
			{8'd132, 8'd97}: color_data = 12'h333;
			{8'd132, 8'd98}: color_data = 12'h333;
			{8'd132, 8'd99}: color_data = 12'h333;
			{8'd132, 8'd100}: color_data = 12'h333;
			{8'd132, 8'd101}: color_data = 12'h333;
			{8'd132, 8'd102}: color_data = 12'h333;
			{8'd132, 8'd103}: color_data = 12'h333;
			{8'd132, 8'd104}: color_data = 12'h333;
			{8'd132, 8'd105}: color_data = 12'h333;
			{8'd132, 8'd106}: color_data = 12'h333;
			{8'd132, 8'd107}: color_data = 12'h333;
			{8'd132, 8'd108}: color_data = 12'h222;
			{8'd132, 8'd109}: color_data = 12'h222;
			{8'd132, 8'd110}: color_data = 12'h222;
			{8'd132, 8'd111}: color_data = 12'h222;
			{8'd132, 8'd112}: color_data = 12'h222;
			{8'd132, 8'd113}: color_data = 12'h222;
			{8'd132, 8'd114}: color_data = 12'h222;
			{8'd132, 8'd115}: color_data = 12'h222;
			{8'd132, 8'd116}: color_data = 12'h222;
			{8'd132, 8'd117}: color_data = 12'h222;
			{8'd132, 8'd118}: color_data = 12'h222;
			{8'd132, 8'd119}: color_data = 12'h222;
			{8'd132, 8'd120}: color_data = 12'h222;
			{8'd132, 8'd121}: color_data = 12'h111;
			{8'd132, 8'd122}: color_data = 12'h111;
			{8'd132, 8'd123}: color_data = 12'h566;
			{8'd132, 8'd124}: color_data = 12'hddd;
			{8'd132, 8'd125}: color_data = 12'h777;
			{8'd132, 8'd126}: color_data = 12'h544;
			{8'd132, 8'd127}: color_data = 12'h421;
			{8'd132, 8'd128}: color_data = 12'h521;
			{8'd132, 8'd129}: color_data = 12'h321;
			{8'd132, 8'd130}: color_data = 12'h999;
			{8'd132, 8'd131}: color_data = 12'hfff;
			{8'd132, 8'd132}: color_data = 12'hfff;
			{8'd132, 8'd133}: color_data = 12'hfff;
			{8'd132, 8'd134}: color_data = 12'hfff;
			{8'd132, 8'd135}: color_data = 12'hfff;
			{8'd132, 8'd136}: color_data = 12'hfff;
			{8'd132, 8'd137}: color_data = 12'hfff;
			{8'd132, 8'd138}: color_data = 12'hfff;
			{8'd132, 8'd139}: color_data = 12'hccc;
			{8'd132, 8'd140}: color_data = 12'h999;
			{8'd133, 8'd18}: color_data = 12'h888;
			{8'd133, 8'd19}: color_data = 12'ha99;
			{8'd133, 8'd20}: color_data = 12'h999;
			{8'd133, 8'd21}: color_data = 12'h999;
			{8'd133, 8'd22}: color_data = 12'h999;
			{8'd133, 8'd23}: color_data = 12'h999;
			{8'd133, 8'd24}: color_data = 12'h999;
			{8'd133, 8'd25}: color_data = 12'h999;
			{8'd133, 8'd26}: color_data = 12'h999;
			{8'd133, 8'd27}: color_data = 12'h999;
			{8'd133, 8'd28}: color_data = 12'h999;
			{8'd133, 8'd29}: color_data = 12'h999;
			{8'd133, 8'd30}: color_data = 12'h999;
			{8'd133, 8'd31}: color_data = 12'h999;
			{8'd133, 8'd32}: color_data = 12'h888;
			{8'd133, 8'd33}: color_data = 12'h777;
			{8'd133, 8'd34}: color_data = 12'h578;
			{8'd133, 8'd35}: color_data = 12'hf00;
			{8'd133, 8'd36}: color_data = 12'hd31;
			{8'd133, 8'd37}: color_data = 12'he41;
			{8'd133, 8'd38}: color_data = 12'he41;
			{8'd133, 8'd39}: color_data = 12'he51;
			{8'd133, 8'd40}: color_data = 12'he51;
			{8'd133, 8'd41}: color_data = 12'he51;
			{8'd133, 8'd42}: color_data = 12'he61;
			{8'd133, 8'd43}: color_data = 12'he61;
			{8'd133, 8'd44}: color_data = 12'he71;
			{8'd133, 8'd45}: color_data = 12'he71;
			{8'd133, 8'd46}: color_data = 12'he71;
			{8'd133, 8'd47}: color_data = 12'he80;
			{8'd133, 8'd48}: color_data = 12'he80;
			{8'd133, 8'd49}: color_data = 12'he80;
			{8'd133, 8'd50}: color_data = 12'hc70;
			{8'd133, 8'd51}: color_data = 12'hc70;
			{8'd133, 8'd53}: color_data = 12'h555;
			{8'd133, 8'd54}: color_data = 12'h666;
			{8'd133, 8'd55}: color_data = 12'h777;
			{8'd133, 8'd56}: color_data = 12'h666;
			{8'd133, 8'd57}: color_data = 12'h666;
			{8'd133, 8'd58}: color_data = 12'h666;
			{8'd133, 8'd59}: color_data = 12'h666;
			{8'd133, 8'd60}: color_data = 12'h666;
			{8'd133, 8'd61}: color_data = 12'h666;
			{8'd133, 8'd62}: color_data = 12'h666;
			{8'd133, 8'd63}: color_data = 12'h666;
			{8'd133, 8'd64}: color_data = 12'h666;
			{8'd133, 8'd65}: color_data = 12'h666;
			{8'd133, 8'd66}: color_data = 12'h666;
			{8'd133, 8'd67}: color_data = 12'h666;
			{8'd133, 8'd68}: color_data = 12'h666;
			{8'd133, 8'd69}: color_data = 12'h555;
			{8'd133, 8'd70}: color_data = 12'h555;
			{8'd133, 8'd71}: color_data = 12'h555;
			{8'd133, 8'd72}: color_data = 12'h555;
			{8'd133, 8'd73}: color_data = 12'h555;
			{8'd133, 8'd74}: color_data = 12'h555;
			{8'd133, 8'd75}: color_data = 12'h555;
			{8'd133, 8'd76}: color_data = 12'h555;
			{8'd133, 8'd77}: color_data = 12'h555;
			{8'd133, 8'd78}: color_data = 12'h555;
			{8'd133, 8'd79}: color_data = 12'h555;
			{8'd133, 8'd80}: color_data = 12'h555;
			{8'd133, 8'd81}: color_data = 12'h444;
			{8'd133, 8'd82}: color_data = 12'h444;
			{8'd133, 8'd83}: color_data = 12'h444;
			{8'd133, 8'd84}: color_data = 12'h444;
			{8'd133, 8'd85}: color_data = 12'h444;
			{8'd133, 8'd86}: color_data = 12'h444;
			{8'd133, 8'd87}: color_data = 12'h444;
			{8'd133, 8'd88}: color_data = 12'h444;
			{8'd133, 8'd89}: color_data = 12'h444;
			{8'd133, 8'd90}: color_data = 12'h444;
			{8'd133, 8'd91}: color_data = 12'h444;
			{8'd133, 8'd92}: color_data = 12'h444;
			{8'd133, 8'd93}: color_data = 12'h444;
			{8'd133, 8'd94}: color_data = 12'h333;
			{8'd133, 8'd95}: color_data = 12'h333;
			{8'd133, 8'd96}: color_data = 12'h333;
			{8'd133, 8'd97}: color_data = 12'h333;
			{8'd133, 8'd98}: color_data = 12'h333;
			{8'd133, 8'd99}: color_data = 12'h333;
			{8'd133, 8'd100}: color_data = 12'h333;
			{8'd133, 8'd101}: color_data = 12'h333;
			{8'd133, 8'd102}: color_data = 12'h333;
			{8'd133, 8'd103}: color_data = 12'h333;
			{8'd133, 8'd104}: color_data = 12'h333;
			{8'd133, 8'd105}: color_data = 12'h333;
			{8'd133, 8'd106}: color_data = 12'h333;
			{8'd133, 8'd107}: color_data = 12'h333;
			{8'd133, 8'd108}: color_data = 12'h222;
			{8'd133, 8'd109}: color_data = 12'h222;
			{8'd133, 8'd110}: color_data = 12'h222;
			{8'd133, 8'd111}: color_data = 12'h222;
			{8'd133, 8'd112}: color_data = 12'h222;
			{8'd133, 8'd113}: color_data = 12'h222;
			{8'd133, 8'd114}: color_data = 12'h222;
			{8'd133, 8'd115}: color_data = 12'h222;
			{8'd133, 8'd116}: color_data = 12'h222;
			{8'd133, 8'd117}: color_data = 12'h222;
			{8'd133, 8'd118}: color_data = 12'h222;
			{8'd133, 8'd119}: color_data = 12'h222;
			{8'd133, 8'd120}: color_data = 12'h222;
			{8'd133, 8'd121}: color_data = 12'h111;
			{8'd133, 8'd122}: color_data = 12'h111;
			{8'd133, 8'd123}: color_data = 12'h444;
			{8'd133, 8'd124}: color_data = 12'hddd;
			{8'd133, 8'd125}: color_data = 12'hfff;
			{8'd133, 8'd126}: color_data = 12'hccc;
			{8'd133, 8'd127}: color_data = 12'h888;
			{8'd133, 8'd128}: color_data = 12'h888;
			{8'd133, 8'd129}: color_data = 12'haaa;
			{8'd133, 8'd130}: color_data = 12'hfff;
			{8'd133, 8'd131}: color_data = 12'hfff;
			{8'd133, 8'd132}: color_data = 12'hfff;
			{8'd133, 8'd133}: color_data = 12'hfff;
			{8'd133, 8'd134}: color_data = 12'hfff;
			{8'd133, 8'd135}: color_data = 12'hfff;
			{8'd133, 8'd136}: color_data = 12'hfff;
			{8'd133, 8'd137}: color_data = 12'hfff;
			{8'd133, 8'd138}: color_data = 12'hfff;
			{8'd133, 8'd139}: color_data = 12'hbbb;
			{8'd133, 8'd140}: color_data = 12'h777;
			{8'd134, 8'd24}: color_data = 12'h999;
			{8'd134, 8'd25}: color_data = 12'h999;
			{8'd134, 8'd26}: color_data = 12'h999;
			{8'd134, 8'd27}: color_data = 12'h999;
			{8'd134, 8'd28}: color_data = 12'h888;
			{8'd134, 8'd29}: color_data = 12'h888;
			{8'd134, 8'd30}: color_data = 12'h888;
			{8'd134, 8'd31}: color_data = 12'h888;
			{8'd134, 8'd32}: color_data = 12'h888;
			{8'd134, 8'd34}: color_data = 12'hc11;
			{8'd134, 8'd35}: color_data = 12'hd21;
			{8'd134, 8'd36}: color_data = 12'hd31;
			{8'd134, 8'd37}: color_data = 12'he41;
			{8'd134, 8'd38}: color_data = 12'he41;
			{8'd134, 8'd39}: color_data = 12'he51;
			{8'd134, 8'd40}: color_data = 12'he51;
			{8'd134, 8'd41}: color_data = 12'he61;
			{8'd134, 8'd42}: color_data = 12'he61;
			{8'd134, 8'd43}: color_data = 12'he61;
			{8'd134, 8'd44}: color_data = 12'he71;
			{8'd134, 8'd45}: color_data = 12'he71;
			{8'd134, 8'd46}: color_data = 12'he71;
			{8'd134, 8'd47}: color_data = 12'he80;
			{8'd134, 8'd48}: color_data = 12'he80;
			{8'd134, 8'd49}: color_data = 12'he80;
			{8'd134, 8'd50}: color_data = 12'he90;
			{8'd134, 8'd51}: color_data = 12'hd80;
			{8'd134, 8'd52}: color_data = 12'hd80;
			{8'd134, 8'd54}: color_data = 12'h666;
			{8'd134, 8'd55}: color_data = 12'h666;
			{8'd134, 8'd56}: color_data = 12'h777;
			{8'd134, 8'd57}: color_data = 12'h666;
			{8'd134, 8'd58}: color_data = 12'h666;
			{8'd134, 8'd59}: color_data = 12'h666;
			{8'd134, 8'd60}: color_data = 12'h666;
			{8'd134, 8'd61}: color_data = 12'h666;
			{8'd134, 8'd62}: color_data = 12'h666;
			{8'd134, 8'd63}: color_data = 12'h666;
			{8'd134, 8'd64}: color_data = 12'h666;
			{8'd134, 8'd65}: color_data = 12'h666;
			{8'd134, 8'd66}: color_data = 12'h666;
			{8'd134, 8'd67}: color_data = 12'h666;
			{8'd134, 8'd68}: color_data = 12'h666;
			{8'd134, 8'd69}: color_data = 12'h555;
			{8'd134, 8'd70}: color_data = 12'h555;
			{8'd134, 8'd71}: color_data = 12'h555;
			{8'd134, 8'd72}: color_data = 12'h555;
			{8'd134, 8'd73}: color_data = 12'h555;
			{8'd134, 8'd74}: color_data = 12'h555;
			{8'd134, 8'd75}: color_data = 12'h555;
			{8'd134, 8'd76}: color_data = 12'h555;
			{8'd134, 8'd77}: color_data = 12'h555;
			{8'd134, 8'd78}: color_data = 12'h555;
			{8'd134, 8'd79}: color_data = 12'h555;
			{8'd134, 8'd80}: color_data = 12'h555;
			{8'd134, 8'd81}: color_data = 12'h444;
			{8'd134, 8'd82}: color_data = 12'h444;
			{8'd134, 8'd83}: color_data = 12'h444;
			{8'd134, 8'd84}: color_data = 12'h444;
			{8'd134, 8'd85}: color_data = 12'h444;
			{8'd134, 8'd86}: color_data = 12'h444;
			{8'd134, 8'd87}: color_data = 12'h444;
			{8'd134, 8'd88}: color_data = 12'h444;
			{8'd134, 8'd89}: color_data = 12'h444;
			{8'd134, 8'd90}: color_data = 12'h444;
			{8'd134, 8'd91}: color_data = 12'h444;
			{8'd134, 8'd92}: color_data = 12'h444;
			{8'd134, 8'd93}: color_data = 12'h444;
			{8'd134, 8'd94}: color_data = 12'h333;
			{8'd134, 8'd95}: color_data = 12'h333;
			{8'd134, 8'd96}: color_data = 12'h333;
			{8'd134, 8'd97}: color_data = 12'h333;
			{8'd134, 8'd98}: color_data = 12'h333;
			{8'd134, 8'd99}: color_data = 12'h333;
			{8'd134, 8'd100}: color_data = 12'h333;
			{8'd134, 8'd101}: color_data = 12'h333;
			{8'd134, 8'd102}: color_data = 12'h333;
			{8'd134, 8'd103}: color_data = 12'h333;
			{8'd134, 8'd104}: color_data = 12'h333;
			{8'd134, 8'd105}: color_data = 12'h333;
			{8'd134, 8'd106}: color_data = 12'h333;
			{8'd134, 8'd107}: color_data = 12'h222;
			{8'd134, 8'd108}: color_data = 12'h222;
			{8'd134, 8'd109}: color_data = 12'h222;
			{8'd134, 8'd110}: color_data = 12'h222;
			{8'd134, 8'd111}: color_data = 12'h222;
			{8'd134, 8'd112}: color_data = 12'h222;
			{8'd134, 8'd113}: color_data = 12'h222;
			{8'd134, 8'd114}: color_data = 12'h222;
			{8'd134, 8'd115}: color_data = 12'h222;
			{8'd134, 8'd116}: color_data = 12'h222;
			{8'd134, 8'd117}: color_data = 12'h222;
			{8'd134, 8'd118}: color_data = 12'h222;
			{8'd134, 8'd119}: color_data = 12'h222;
			{8'd134, 8'd120}: color_data = 12'h222;
			{8'd134, 8'd121}: color_data = 12'h111;
			{8'd134, 8'd122}: color_data = 12'h111;
			{8'd134, 8'd123}: color_data = 12'h333;
			{8'd134, 8'd124}: color_data = 12'hccc;
			{8'd134, 8'd125}: color_data = 12'hfff;
			{8'd134, 8'd126}: color_data = 12'hfff;
			{8'd134, 8'd127}: color_data = 12'hfff;
			{8'd134, 8'd128}: color_data = 12'hfff;
			{8'd134, 8'd129}: color_data = 12'hfff;
			{8'd134, 8'd130}: color_data = 12'hfff;
			{8'd134, 8'd131}: color_data = 12'hfff;
			{8'd134, 8'd132}: color_data = 12'hfff;
			{8'd134, 8'd133}: color_data = 12'hfff;
			{8'd134, 8'd134}: color_data = 12'hfff;
			{8'd134, 8'd135}: color_data = 12'hfff;
			{8'd134, 8'd136}: color_data = 12'hfff;
			{8'd134, 8'd137}: color_data = 12'hfff;
			{8'd134, 8'd138}: color_data = 12'hfff;
			{8'd134, 8'd139}: color_data = 12'haaa;
			{8'd134, 8'd140}: color_data = 12'h666;
			{8'd135, 8'd28}: color_data = 12'h777;
			{8'd135, 8'd29}: color_data = 12'h777;
			{8'd135, 8'd30}: color_data = 12'h888;
			{8'd135, 8'd31}: color_data = 12'h888;
			{8'd135, 8'd32}: color_data = 12'h5aa;
			{8'd135, 8'd33}: color_data = 12'hb11;
			{8'd135, 8'd34}: color_data = 12'hc21;
			{8'd135, 8'd35}: color_data = 12'he21;
			{8'd135, 8'd36}: color_data = 12'hd31;
			{8'd135, 8'd37}: color_data = 12'hd41;
			{8'd135, 8'd38}: color_data = 12'he41;
			{8'd135, 8'd39}: color_data = 12'hd41;
			{8'd135, 8'd40}: color_data = 12'hd41;
			{8'd135, 8'd41}: color_data = 12'hd51;
			{8'd135, 8'd42}: color_data = 12'he61;
			{8'd135, 8'd43}: color_data = 12'he61;
			{8'd135, 8'd44}: color_data = 12'hd61;
			{8'd135, 8'd45}: color_data = 12'hd71;
			{8'd135, 8'd46}: color_data = 12'he71;
			{8'd135, 8'd47}: color_data = 12'he80;
			{8'd135, 8'd48}: color_data = 12'he80;
			{8'd135, 8'd49}: color_data = 12'he80;
			{8'd135, 8'd50}: color_data = 12'he90;
			{8'd135, 8'd51}: color_data = 12'he90;
			{8'd135, 8'd52}: color_data = 12'hd90;
			{8'd135, 8'd53}: color_data = 12'hfa0;
			{8'd135, 8'd54}: color_data = 12'h667;
			{8'd135, 8'd55}: color_data = 12'h777;
			{8'd135, 8'd56}: color_data = 12'h777;
			{8'd135, 8'd57}: color_data = 12'h666;
			{8'd135, 8'd58}: color_data = 12'h666;
			{8'd135, 8'd59}: color_data = 12'h666;
			{8'd135, 8'd60}: color_data = 12'h666;
			{8'd135, 8'd61}: color_data = 12'h666;
			{8'd135, 8'd62}: color_data = 12'h666;
			{8'd135, 8'd63}: color_data = 12'h666;
			{8'd135, 8'd64}: color_data = 12'h666;
			{8'd135, 8'd65}: color_data = 12'h666;
			{8'd135, 8'd66}: color_data = 12'h666;
			{8'd135, 8'd67}: color_data = 12'h666;
			{8'd135, 8'd68}: color_data = 12'h555;
			{8'd135, 8'd69}: color_data = 12'h555;
			{8'd135, 8'd70}: color_data = 12'h555;
			{8'd135, 8'd71}: color_data = 12'h555;
			{8'd135, 8'd72}: color_data = 12'h555;
			{8'd135, 8'd73}: color_data = 12'h555;
			{8'd135, 8'd74}: color_data = 12'h555;
			{8'd135, 8'd75}: color_data = 12'h555;
			{8'd135, 8'd76}: color_data = 12'h555;
			{8'd135, 8'd77}: color_data = 12'h555;
			{8'd135, 8'd78}: color_data = 12'h555;
			{8'd135, 8'd79}: color_data = 12'h555;
			{8'd135, 8'd80}: color_data = 12'h555;
			{8'd135, 8'd81}: color_data = 12'h444;
			{8'd135, 8'd82}: color_data = 12'h444;
			{8'd135, 8'd83}: color_data = 12'h444;
			{8'd135, 8'd84}: color_data = 12'h444;
			{8'd135, 8'd85}: color_data = 12'h444;
			{8'd135, 8'd86}: color_data = 12'h444;
			{8'd135, 8'd87}: color_data = 12'h444;
			{8'd135, 8'd88}: color_data = 12'h444;
			{8'd135, 8'd89}: color_data = 12'h444;
			{8'd135, 8'd90}: color_data = 12'h444;
			{8'd135, 8'd91}: color_data = 12'h444;
			{8'd135, 8'd92}: color_data = 12'h444;
			{8'd135, 8'd93}: color_data = 12'h444;
			{8'd135, 8'd94}: color_data = 12'h333;
			{8'd135, 8'd95}: color_data = 12'h333;
			{8'd135, 8'd96}: color_data = 12'h333;
			{8'd135, 8'd97}: color_data = 12'h333;
			{8'd135, 8'd98}: color_data = 12'h333;
			{8'd135, 8'd99}: color_data = 12'h333;
			{8'd135, 8'd100}: color_data = 12'h333;
			{8'd135, 8'd101}: color_data = 12'h333;
			{8'd135, 8'd102}: color_data = 12'h333;
			{8'd135, 8'd103}: color_data = 12'h333;
			{8'd135, 8'd104}: color_data = 12'h333;
			{8'd135, 8'd105}: color_data = 12'h333;
			{8'd135, 8'd106}: color_data = 12'h333;
			{8'd135, 8'd107}: color_data = 12'h222;
			{8'd135, 8'd108}: color_data = 12'h222;
			{8'd135, 8'd109}: color_data = 12'h222;
			{8'd135, 8'd110}: color_data = 12'h222;
			{8'd135, 8'd111}: color_data = 12'h222;
			{8'd135, 8'd112}: color_data = 12'h222;
			{8'd135, 8'd113}: color_data = 12'h222;
			{8'd135, 8'd114}: color_data = 12'h222;
			{8'd135, 8'd115}: color_data = 12'h222;
			{8'd135, 8'd116}: color_data = 12'h222;
			{8'd135, 8'd117}: color_data = 12'h222;
			{8'd135, 8'd118}: color_data = 12'h222;
			{8'd135, 8'd119}: color_data = 12'h222;
			{8'd135, 8'd120}: color_data = 12'h222;
			{8'd135, 8'd121}: color_data = 12'h111;
			{8'd135, 8'd122}: color_data = 12'h111;
			{8'd135, 8'd123}: color_data = 12'h222;
			{8'd135, 8'd124}: color_data = 12'haaa;
			{8'd135, 8'd125}: color_data = 12'hfff;
			{8'd135, 8'd126}: color_data = 12'hfff;
			{8'd135, 8'd127}: color_data = 12'hfff;
			{8'd135, 8'd128}: color_data = 12'hfff;
			{8'd135, 8'd129}: color_data = 12'hfff;
			{8'd135, 8'd130}: color_data = 12'hfff;
			{8'd135, 8'd131}: color_data = 12'hfff;
			{8'd135, 8'd132}: color_data = 12'hfff;
			{8'd135, 8'd133}: color_data = 12'hfff;
			{8'd135, 8'd134}: color_data = 12'hfff;
			{8'd135, 8'd135}: color_data = 12'hfff;
			{8'd135, 8'd136}: color_data = 12'hfff;
			{8'd135, 8'd137}: color_data = 12'hfff;
			{8'd135, 8'd138}: color_data = 12'heee;
			{8'd135, 8'd139}: color_data = 12'h999;
			{8'd135, 8'd140}: color_data = 12'h555;
			{8'd136, 8'd32}: color_data = 12'ha01;
			{8'd136, 8'd33}: color_data = 12'hc11;
			{8'd136, 8'd34}: color_data = 12'he21;
			{8'd136, 8'd35}: color_data = 12'hd21;
			{8'd136, 8'd36}: color_data = 12'hd31;
			{8'd136, 8'd37}: color_data = 12'hd41;
			{8'd136, 8'd38}: color_data = 12'he41;
			{8'd136, 8'd39}: color_data = 12'hb30;
			{8'd136, 8'd40}: color_data = 12'h930;
			{8'd136, 8'd41}: color_data = 12'hc41;
			{8'd136, 8'd42}: color_data = 12'hd61;
			{8'd136, 8'd43}: color_data = 12'hc61;
			{8'd136, 8'd44}: color_data = 12'ha51;
			{8'd136, 8'd45}: color_data = 12'hb61;
			{8'd136, 8'd46}: color_data = 12'hd71;
			{8'd136, 8'd47}: color_data = 12'he80;
			{8'd136, 8'd48}: color_data = 12'he80;
			{8'd136, 8'd49}: color_data = 12'he80;
			{8'd136, 8'd50}: color_data = 12'he90;
			{8'd136, 8'd51}: color_data = 12'he90;
			{8'd136, 8'd52}: color_data = 12'hd90;
			{8'd136, 8'd53}: color_data = 12'hd80;
			{8'd136, 8'd54}: color_data = 12'h667;
			{8'd136, 8'd55}: color_data = 12'h777;
			{8'd136, 8'd56}: color_data = 12'h777;
			{8'd136, 8'd57}: color_data = 12'h666;
			{8'd136, 8'd58}: color_data = 12'h666;
			{8'd136, 8'd59}: color_data = 12'h666;
			{8'd136, 8'd60}: color_data = 12'h666;
			{8'd136, 8'd61}: color_data = 12'h666;
			{8'd136, 8'd62}: color_data = 12'h666;
			{8'd136, 8'd63}: color_data = 12'h666;
			{8'd136, 8'd64}: color_data = 12'h666;
			{8'd136, 8'd65}: color_data = 12'h666;
			{8'd136, 8'd66}: color_data = 12'h666;
			{8'd136, 8'd67}: color_data = 12'h666;
			{8'd136, 8'd68}: color_data = 12'h555;
			{8'd136, 8'd69}: color_data = 12'h555;
			{8'd136, 8'd70}: color_data = 12'h555;
			{8'd136, 8'd71}: color_data = 12'h555;
			{8'd136, 8'd72}: color_data = 12'h555;
			{8'd136, 8'd73}: color_data = 12'h555;
			{8'd136, 8'd74}: color_data = 12'h555;
			{8'd136, 8'd75}: color_data = 12'h555;
			{8'd136, 8'd76}: color_data = 12'h555;
			{8'd136, 8'd77}: color_data = 12'h555;
			{8'd136, 8'd78}: color_data = 12'h555;
			{8'd136, 8'd79}: color_data = 12'h555;
			{8'd136, 8'd80}: color_data = 12'h555;
			{8'd136, 8'd81}: color_data = 12'h444;
			{8'd136, 8'd82}: color_data = 12'h444;
			{8'd136, 8'd83}: color_data = 12'h444;
			{8'd136, 8'd84}: color_data = 12'h444;
			{8'd136, 8'd85}: color_data = 12'h444;
			{8'd136, 8'd86}: color_data = 12'h444;
			{8'd136, 8'd87}: color_data = 12'h444;
			{8'd136, 8'd88}: color_data = 12'h444;
			{8'd136, 8'd89}: color_data = 12'h444;
			{8'd136, 8'd90}: color_data = 12'h444;
			{8'd136, 8'd91}: color_data = 12'h444;
			{8'd136, 8'd92}: color_data = 12'h444;
			{8'd136, 8'd93}: color_data = 12'h444;
			{8'd136, 8'd94}: color_data = 12'h333;
			{8'd136, 8'd95}: color_data = 12'h333;
			{8'd136, 8'd96}: color_data = 12'h333;
			{8'd136, 8'd97}: color_data = 12'h333;
			{8'd136, 8'd98}: color_data = 12'h333;
			{8'd136, 8'd99}: color_data = 12'h333;
			{8'd136, 8'd100}: color_data = 12'h333;
			{8'd136, 8'd101}: color_data = 12'h333;
			{8'd136, 8'd102}: color_data = 12'h333;
			{8'd136, 8'd103}: color_data = 12'h333;
			{8'd136, 8'd104}: color_data = 12'h333;
			{8'd136, 8'd105}: color_data = 12'h333;
			{8'd136, 8'd106}: color_data = 12'h333;
			{8'd136, 8'd107}: color_data = 12'h222;
			{8'd136, 8'd108}: color_data = 12'h222;
			{8'd136, 8'd109}: color_data = 12'h222;
			{8'd136, 8'd110}: color_data = 12'h222;
			{8'd136, 8'd111}: color_data = 12'h222;
			{8'd136, 8'd112}: color_data = 12'h222;
			{8'd136, 8'd113}: color_data = 12'h222;
			{8'd136, 8'd114}: color_data = 12'h222;
			{8'd136, 8'd115}: color_data = 12'h222;
			{8'd136, 8'd116}: color_data = 12'h222;
			{8'd136, 8'd117}: color_data = 12'h222;
			{8'd136, 8'd118}: color_data = 12'h222;
			{8'd136, 8'd119}: color_data = 12'h222;
			{8'd136, 8'd120}: color_data = 12'h222;
			{8'd136, 8'd121}: color_data = 12'h111;
			{8'd136, 8'd122}: color_data = 12'h111;
			{8'd136, 8'd123}: color_data = 12'h111;
			{8'd136, 8'd124}: color_data = 12'h888;
			{8'd136, 8'd125}: color_data = 12'hfff;
			{8'd136, 8'd126}: color_data = 12'hfff;
			{8'd136, 8'd127}: color_data = 12'hfff;
			{8'd136, 8'd128}: color_data = 12'hfff;
			{8'd136, 8'd129}: color_data = 12'hfff;
			{8'd136, 8'd130}: color_data = 12'hfff;
			{8'd136, 8'd131}: color_data = 12'hfff;
			{8'd136, 8'd132}: color_data = 12'hfff;
			{8'd136, 8'd133}: color_data = 12'hfff;
			{8'd136, 8'd134}: color_data = 12'hfff;
			{8'd136, 8'd135}: color_data = 12'hfff;
			{8'd136, 8'd136}: color_data = 12'hfff;
			{8'd136, 8'd137}: color_data = 12'hfff;
			{8'd136, 8'd138}: color_data = 12'heee;
			{8'd136, 8'd139}: color_data = 12'h999;
			{8'd136, 8'd140}: color_data = 12'h555;
			{8'd137, 8'd32}: color_data = 12'hb11;
			{8'd137, 8'd33}: color_data = 12'hd11;
			{8'd137, 8'd34}: color_data = 12'hd21;
			{8'd137, 8'd35}: color_data = 12'hd21;
			{8'd137, 8'd36}: color_data = 12'hd31;
			{8'd137, 8'd37}: color_data = 12'he41;
			{8'd137, 8'd38}: color_data = 12'hc41;
			{8'd137, 8'd39}: color_data = 12'h930;
			{8'd137, 8'd45}: color_data = 12'h840;
			{8'd137, 8'd46}: color_data = 12'ha50;
			{8'd137, 8'd47}: color_data = 12'hd70;
			{8'd137, 8'd48}: color_data = 12'he80;
			{8'd137, 8'd49}: color_data = 12'he80;
			{8'd137, 8'd50}: color_data = 12'he90;
			{8'd137, 8'd51}: color_data = 12'he90;
			{8'd137, 8'd52}: color_data = 12'hd90;
			{8'd137, 8'd53}: color_data = 12'hd80;
			{8'd137, 8'd54}: color_data = 12'h667;
			{8'd137, 8'd55}: color_data = 12'h666;
			{8'd137, 8'd56}: color_data = 12'h666;
			{8'd137, 8'd57}: color_data = 12'h666;
			{8'd137, 8'd58}: color_data = 12'h666;
			{8'd137, 8'd59}: color_data = 12'h666;
			{8'd137, 8'd60}: color_data = 12'h666;
			{8'd137, 8'd61}: color_data = 12'h666;
			{8'd137, 8'd62}: color_data = 12'h666;
			{8'd137, 8'd63}: color_data = 12'h666;
			{8'd137, 8'd64}: color_data = 12'h666;
			{8'd137, 8'd65}: color_data = 12'h666;
			{8'd137, 8'd66}: color_data = 12'h666;
			{8'd137, 8'd67}: color_data = 12'h666;
			{8'd137, 8'd68}: color_data = 12'h555;
			{8'd137, 8'd69}: color_data = 12'h555;
			{8'd137, 8'd70}: color_data = 12'h555;
			{8'd137, 8'd71}: color_data = 12'h555;
			{8'd137, 8'd72}: color_data = 12'h555;
			{8'd137, 8'd73}: color_data = 12'h555;
			{8'd137, 8'd74}: color_data = 12'h555;
			{8'd137, 8'd75}: color_data = 12'h555;
			{8'd137, 8'd76}: color_data = 12'h555;
			{8'd137, 8'd77}: color_data = 12'h555;
			{8'd137, 8'd78}: color_data = 12'h555;
			{8'd137, 8'd79}: color_data = 12'h555;
			{8'd137, 8'd80}: color_data = 12'h555;
			{8'd137, 8'd81}: color_data = 12'h444;
			{8'd137, 8'd82}: color_data = 12'h444;
			{8'd137, 8'd83}: color_data = 12'h444;
			{8'd137, 8'd84}: color_data = 12'h444;
			{8'd137, 8'd85}: color_data = 12'h444;
			{8'd137, 8'd86}: color_data = 12'h444;
			{8'd137, 8'd87}: color_data = 12'h444;
			{8'd137, 8'd88}: color_data = 12'h444;
			{8'd137, 8'd89}: color_data = 12'h444;
			{8'd137, 8'd90}: color_data = 12'h444;
			{8'd137, 8'd91}: color_data = 12'h444;
			{8'd137, 8'd92}: color_data = 12'h444;
			{8'd137, 8'd93}: color_data = 12'h444;
			{8'd137, 8'd94}: color_data = 12'h333;
			{8'd137, 8'd95}: color_data = 12'h333;
			{8'd137, 8'd96}: color_data = 12'h333;
			{8'd137, 8'd97}: color_data = 12'h333;
			{8'd137, 8'd98}: color_data = 12'h333;
			{8'd137, 8'd99}: color_data = 12'h333;
			{8'd137, 8'd100}: color_data = 12'h333;
			{8'd137, 8'd101}: color_data = 12'h333;
			{8'd137, 8'd102}: color_data = 12'h333;
			{8'd137, 8'd103}: color_data = 12'h333;
			{8'd137, 8'd104}: color_data = 12'h333;
			{8'd137, 8'd105}: color_data = 12'h333;
			{8'd137, 8'd106}: color_data = 12'h333;
			{8'd137, 8'd107}: color_data = 12'h222;
			{8'd137, 8'd108}: color_data = 12'h222;
			{8'd137, 8'd109}: color_data = 12'h222;
			{8'd137, 8'd110}: color_data = 12'h222;
			{8'd137, 8'd111}: color_data = 12'h222;
			{8'd137, 8'd112}: color_data = 12'h222;
			{8'd137, 8'd113}: color_data = 12'h222;
			{8'd137, 8'd114}: color_data = 12'h222;
			{8'd137, 8'd115}: color_data = 12'h222;
			{8'd137, 8'd116}: color_data = 12'h222;
			{8'd137, 8'd117}: color_data = 12'h222;
			{8'd137, 8'd118}: color_data = 12'h222;
			{8'd137, 8'd119}: color_data = 12'h222;
			{8'd137, 8'd120}: color_data = 12'h222;
			{8'd137, 8'd121}: color_data = 12'h111;
			{8'd137, 8'd122}: color_data = 12'h111;
			{8'd137, 8'd123}: color_data = 12'h111;
			{8'd137, 8'd124}: color_data = 12'h666;
			{8'd137, 8'd125}: color_data = 12'heee;
			{8'd137, 8'd126}: color_data = 12'hfff;
			{8'd137, 8'd127}: color_data = 12'hfff;
			{8'd137, 8'd128}: color_data = 12'hfff;
			{8'd137, 8'd129}: color_data = 12'hfff;
			{8'd137, 8'd130}: color_data = 12'hfff;
			{8'd137, 8'd131}: color_data = 12'hfff;
			{8'd137, 8'd132}: color_data = 12'hfff;
			{8'd137, 8'd133}: color_data = 12'hfff;
			{8'd137, 8'd134}: color_data = 12'hfff;
			{8'd137, 8'd135}: color_data = 12'hfff;
			{8'd137, 8'd136}: color_data = 12'hfff;
			{8'd137, 8'd137}: color_data = 12'hfff;
			{8'd137, 8'd138}: color_data = 12'hddd;
			{8'd137, 8'd139}: color_data = 12'h888;
			{8'd137, 8'd140}: color_data = 12'h000;
			{8'd138, 8'd32}: color_data = 12'ha11;
			{8'd138, 8'd33}: color_data = 12'hd11;
			{8'd138, 8'd34}: color_data = 12'hd21;
			{8'd138, 8'd35}: color_data = 12'hd21;
			{8'd138, 8'd36}: color_data = 12'hd31;
			{8'd138, 8'd37}: color_data = 12'hd31;
			{8'd138, 8'd38}: color_data = 12'ha20;
			{8'd138, 8'd46}: color_data = 12'h740;
			{8'd138, 8'd47}: color_data = 12'hb60;
			{8'd138, 8'd48}: color_data = 12'he80;
			{8'd138, 8'd49}: color_data = 12'he80;
			{8'd138, 8'd50}: color_data = 12'he90;
			{8'd138, 8'd51}: color_data = 12'he90;
			{8'd138, 8'd52}: color_data = 12'hd90;
			{8'd138, 8'd53}: color_data = 12'hd80;
			{8'd138, 8'd54}: color_data = 12'h667;
			{8'd138, 8'd55}: color_data = 12'h777;
			{8'd138, 8'd56}: color_data = 12'h777;
			{8'd138, 8'd57}: color_data = 12'h666;
			{8'd138, 8'd58}: color_data = 12'h666;
			{8'd138, 8'd59}: color_data = 12'h666;
			{8'd138, 8'd60}: color_data = 12'h666;
			{8'd138, 8'd61}: color_data = 12'h666;
			{8'd138, 8'd62}: color_data = 12'h666;
			{8'd138, 8'd63}: color_data = 12'h666;
			{8'd138, 8'd64}: color_data = 12'h666;
			{8'd138, 8'd65}: color_data = 12'h666;
			{8'd138, 8'd66}: color_data = 12'h666;
			{8'd138, 8'd67}: color_data = 12'h666;
			{8'd138, 8'd68}: color_data = 12'h555;
			{8'd138, 8'd69}: color_data = 12'h555;
			{8'd138, 8'd70}: color_data = 12'h555;
			{8'd138, 8'd71}: color_data = 12'h555;
			{8'd138, 8'd72}: color_data = 12'h555;
			{8'd138, 8'd73}: color_data = 12'h555;
			{8'd138, 8'd74}: color_data = 12'h555;
			{8'd138, 8'd75}: color_data = 12'h555;
			{8'd138, 8'd76}: color_data = 12'h555;
			{8'd138, 8'd77}: color_data = 12'h555;
			{8'd138, 8'd78}: color_data = 12'h555;
			{8'd138, 8'd79}: color_data = 12'h555;
			{8'd138, 8'd80}: color_data = 12'h555;
			{8'd138, 8'd81}: color_data = 12'h444;
			{8'd138, 8'd82}: color_data = 12'h444;
			{8'd138, 8'd83}: color_data = 12'h444;
			{8'd138, 8'd84}: color_data = 12'h444;
			{8'd138, 8'd85}: color_data = 12'h444;
			{8'd138, 8'd86}: color_data = 12'h444;
			{8'd138, 8'd87}: color_data = 12'h444;
			{8'd138, 8'd88}: color_data = 12'h444;
			{8'd138, 8'd89}: color_data = 12'h444;
			{8'd138, 8'd90}: color_data = 12'h444;
			{8'd138, 8'd91}: color_data = 12'h444;
			{8'd138, 8'd92}: color_data = 12'h444;
			{8'd138, 8'd93}: color_data = 12'h444;
			{8'd138, 8'd94}: color_data = 12'h333;
			{8'd138, 8'd95}: color_data = 12'h333;
			{8'd138, 8'd96}: color_data = 12'h333;
			{8'd138, 8'd97}: color_data = 12'h333;
			{8'd138, 8'd98}: color_data = 12'h333;
			{8'd138, 8'd99}: color_data = 12'h333;
			{8'd138, 8'd100}: color_data = 12'h333;
			{8'd138, 8'd101}: color_data = 12'h333;
			{8'd138, 8'd102}: color_data = 12'h333;
			{8'd138, 8'd103}: color_data = 12'h333;
			{8'd138, 8'd104}: color_data = 12'h333;
			{8'd138, 8'd105}: color_data = 12'h333;
			{8'd138, 8'd106}: color_data = 12'h333;
			{8'd138, 8'd107}: color_data = 12'h222;
			{8'd138, 8'd108}: color_data = 12'h222;
			{8'd138, 8'd109}: color_data = 12'h222;
			{8'd138, 8'd110}: color_data = 12'h222;
			{8'd138, 8'd111}: color_data = 12'h222;
			{8'd138, 8'd112}: color_data = 12'h222;
			{8'd138, 8'd113}: color_data = 12'h222;
			{8'd138, 8'd114}: color_data = 12'h222;
			{8'd138, 8'd115}: color_data = 12'h222;
			{8'd138, 8'd116}: color_data = 12'h222;
			{8'd138, 8'd117}: color_data = 12'h222;
			{8'd138, 8'd118}: color_data = 12'h222;
			{8'd138, 8'd119}: color_data = 12'h222;
			{8'd138, 8'd120}: color_data = 12'h222;
			{8'd138, 8'd121}: color_data = 12'h111;
			{8'd138, 8'd122}: color_data = 12'h111;
			{8'd138, 8'd123}: color_data = 12'h111;
			{8'd138, 8'd124}: color_data = 12'h555;
			{8'd138, 8'd125}: color_data = 12'heee;
			{8'd138, 8'd126}: color_data = 12'hfff;
			{8'd138, 8'd127}: color_data = 12'hfff;
			{8'd138, 8'd128}: color_data = 12'hfff;
			{8'd138, 8'd129}: color_data = 12'hfff;
			{8'd138, 8'd130}: color_data = 12'hfff;
			{8'd138, 8'd131}: color_data = 12'hfff;
			{8'd138, 8'd132}: color_data = 12'hfff;
			{8'd138, 8'd133}: color_data = 12'hfff;
			{8'd138, 8'd134}: color_data = 12'hfff;
			{8'd138, 8'd135}: color_data = 12'hfff;
			{8'd138, 8'd136}: color_data = 12'hfff;
			{8'd138, 8'd137}: color_data = 12'hfff;
			{8'd138, 8'd138}: color_data = 12'hccc;
			{8'd138, 8'd139}: color_data = 12'h777;
			{8'd138, 8'd140}: color_data = 12'h000;
			{8'd139, 8'd32}: color_data = 12'ha11;
			{8'd139, 8'd33}: color_data = 12'hd11;
			{8'd139, 8'd34}: color_data = 12'hd21;
			{8'd139, 8'd35}: color_data = 12'hd21;
			{8'd139, 8'd36}: color_data = 12'hd31;
			{8'd139, 8'd37}: color_data = 12'ha21;
			{8'd139, 8'd38}: color_data = 12'h610;
			{8'd139, 8'd46}: color_data = 12'h950;
			{8'd139, 8'd47}: color_data = 12'hc60;
			{8'd139, 8'd48}: color_data = 12'he80;
			{8'd139, 8'd49}: color_data = 12'he80;
			{8'd139, 8'd50}: color_data = 12'he90;
			{8'd139, 8'd51}: color_data = 12'he90;
			{8'd139, 8'd52}: color_data = 12'hd90;
			{8'd139, 8'd53}: color_data = 12'hc80;
			{8'd139, 8'd54}: color_data = 12'h459;
			{8'd139, 8'd55}: color_data = 12'h666;
			{8'd139, 8'd56}: color_data = 12'h666;
			{8'd139, 8'd57}: color_data = 12'h666;
			{8'd139, 8'd58}: color_data = 12'h666;
			{8'd139, 8'd59}: color_data = 12'h666;
			{8'd139, 8'd60}: color_data = 12'h666;
			{8'd139, 8'd61}: color_data = 12'h666;
			{8'd139, 8'd62}: color_data = 12'h666;
			{8'd139, 8'd63}: color_data = 12'h666;
			{8'd139, 8'd64}: color_data = 12'h666;
			{8'd139, 8'd65}: color_data = 12'h666;
			{8'd139, 8'd66}: color_data = 12'h666;
			{8'd139, 8'd67}: color_data = 12'h666;
			{8'd139, 8'd68}: color_data = 12'h555;
			{8'd139, 8'd69}: color_data = 12'h555;
			{8'd139, 8'd70}: color_data = 12'h555;
			{8'd139, 8'd71}: color_data = 12'h555;
			{8'd139, 8'd72}: color_data = 12'h555;
			{8'd139, 8'd73}: color_data = 12'h555;
			{8'd139, 8'd74}: color_data = 12'h555;
			{8'd139, 8'd75}: color_data = 12'h555;
			{8'd139, 8'd76}: color_data = 12'h555;
			{8'd139, 8'd77}: color_data = 12'h555;
			{8'd139, 8'd78}: color_data = 12'h555;
			{8'd139, 8'd79}: color_data = 12'h555;
			{8'd139, 8'd80}: color_data = 12'h555;
			{8'd139, 8'd81}: color_data = 12'h444;
			{8'd139, 8'd82}: color_data = 12'h444;
			{8'd139, 8'd83}: color_data = 12'h444;
			{8'd139, 8'd84}: color_data = 12'h444;
			{8'd139, 8'd85}: color_data = 12'h444;
			{8'd139, 8'd86}: color_data = 12'h444;
			{8'd139, 8'd87}: color_data = 12'h444;
			{8'd139, 8'd88}: color_data = 12'h444;
			{8'd139, 8'd89}: color_data = 12'h444;
			{8'd139, 8'd90}: color_data = 12'h444;
			{8'd139, 8'd91}: color_data = 12'h444;
			{8'd139, 8'd92}: color_data = 12'h444;
			{8'd139, 8'd93}: color_data = 12'h444;
			{8'd139, 8'd94}: color_data = 12'h333;
			{8'd139, 8'd95}: color_data = 12'h333;
			{8'd139, 8'd96}: color_data = 12'h333;
			{8'd139, 8'd97}: color_data = 12'h333;
			{8'd139, 8'd98}: color_data = 12'h333;
			{8'd139, 8'd99}: color_data = 12'h333;
			{8'd139, 8'd100}: color_data = 12'h333;
			{8'd139, 8'd101}: color_data = 12'h333;
			{8'd139, 8'd102}: color_data = 12'h333;
			{8'd139, 8'd103}: color_data = 12'h333;
			{8'd139, 8'd104}: color_data = 12'h333;
			{8'd139, 8'd105}: color_data = 12'h333;
			{8'd139, 8'd106}: color_data = 12'h333;
			{8'd139, 8'd107}: color_data = 12'h222;
			{8'd139, 8'd108}: color_data = 12'h222;
			{8'd139, 8'd109}: color_data = 12'h222;
			{8'd139, 8'd110}: color_data = 12'h222;
			{8'd139, 8'd111}: color_data = 12'h222;
			{8'd139, 8'd112}: color_data = 12'h222;
			{8'd139, 8'd113}: color_data = 12'h222;
			{8'd139, 8'd114}: color_data = 12'h222;
			{8'd139, 8'd115}: color_data = 12'h222;
			{8'd139, 8'd116}: color_data = 12'h222;
			{8'd139, 8'd117}: color_data = 12'h222;
			{8'd139, 8'd118}: color_data = 12'h222;
			{8'd139, 8'd119}: color_data = 12'h222;
			{8'd139, 8'd120}: color_data = 12'h222;
			{8'd139, 8'd121}: color_data = 12'h111;
			{8'd139, 8'd122}: color_data = 12'h111;
			{8'd139, 8'd123}: color_data = 12'h111;
			{8'd139, 8'd124}: color_data = 12'h333;
			{8'd139, 8'd125}: color_data = 12'hccc;
			{8'd139, 8'd126}: color_data = 12'hfff;
			{8'd139, 8'd127}: color_data = 12'hfff;
			{8'd139, 8'd128}: color_data = 12'hfff;
			{8'd139, 8'd129}: color_data = 12'hfff;
			{8'd139, 8'd130}: color_data = 12'hfff;
			{8'd139, 8'd131}: color_data = 12'hfff;
			{8'd139, 8'd132}: color_data = 12'hfff;
			{8'd139, 8'd133}: color_data = 12'hfff;
			{8'd139, 8'd134}: color_data = 12'hfff;
			{8'd139, 8'd135}: color_data = 12'hfff;
			{8'd139, 8'd136}: color_data = 12'hfff;
			{8'd139, 8'd137}: color_data = 12'hfff;
			{8'd139, 8'd138}: color_data = 12'haaa;
			{8'd139, 8'd139}: color_data = 12'h666;
			{8'd140, 8'd32}: color_data = 12'ha11;
			{8'd140, 8'd33}: color_data = 12'hd11;
			{8'd140, 8'd34}: color_data = 12'hd21;
			{8'd140, 8'd35}: color_data = 12'hd21;
			{8'd140, 8'd36}: color_data = 12'hd31;
			{8'd140, 8'd37}: color_data = 12'ha20;
			{8'd140, 8'd45}: color_data = 12'h951;
			{8'd140, 8'd46}: color_data = 12'hb60;
			{8'd140, 8'd47}: color_data = 12'hd70;
			{8'd140, 8'd48}: color_data = 12'he80;
			{8'd140, 8'd49}: color_data = 12'he80;
			{8'd140, 8'd50}: color_data = 12'he90;
			{8'd140, 8'd51}: color_data = 12'he90;
			{8'd140, 8'd52}: color_data = 12'hd90;
			{8'd140, 8'd53}: color_data = 12'hb80;
			{8'd140, 8'd55}: color_data = 12'h777;
			{8'd140, 8'd56}: color_data = 12'h666;
			{8'd140, 8'd57}: color_data = 12'h777;
			{8'd140, 8'd58}: color_data = 12'h666;
			{8'd140, 8'd59}: color_data = 12'h666;
			{8'd140, 8'd60}: color_data = 12'h666;
			{8'd140, 8'd61}: color_data = 12'h666;
			{8'd140, 8'd62}: color_data = 12'h666;
			{8'd140, 8'd63}: color_data = 12'h666;
			{8'd140, 8'd64}: color_data = 12'h666;
			{8'd140, 8'd65}: color_data = 12'h666;
			{8'd140, 8'd66}: color_data = 12'h666;
			{8'd140, 8'd67}: color_data = 12'h666;
			{8'd140, 8'd68}: color_data = 12'h555;
			{8'd140, 8'd69}: color_data = 12'h555;
			{8'd140, 8'd70}: color_data = 12'h555;
			{8'd140, 8'd71}: color_data = 12'h555;
			{8'd140, 8'd72}: color_data = 12'h555;
			{8'd140, 8'd73}: color_data = 12'h555;
			{8'd140, 8'd74}: color_data = 12'h555;
			{8'd140, 8'd75}: color_data = 12'h555;
			{8'd140, 8'd76}: color_data = 12'h555;
			{8'd140, 8'd77}: color_data = 12'h555;
			{8'd140, 8'd78}: color_data = 12'h555;
			{8'd140, 8'd79}: color_data = 12'h555;
			{8'd140, 8'd80}: color_data = 12'h444;
			{8'd140, 8'd81}: color_data = 12'h444;
			{8'd140, 8'd82}: color_data = 12'h444;
			{8'd140, 8'd83}: color_data = 12'h444;
			{8'd140, 8'd84}: color_data = 12'h444;
			{8'd140, 8'd85}: color_data = 12'h444;
			{8'd140, 8'd86}: color_data = 12'h444;
			{8'd140, 8'd87}: color_data = 12'h444;
			{8'd140, 8'd88}: color_data = 12'h444;
			{8'd140, 8'd89}: color_data = 12'h444;
			{8'd140, 8'd90}: color_data = 12'h444;
			{8'd140, 8'd91}: color_data = 12'h444;
			{8'd140, 8'd92}: color_data = 12'h444;
			{8'd140, 8'd93}: color_data = 12'h333;
			{8'd140, 8'd94}: color_data = 12'h333;
			{8'd140, 8'd95}: color_data = 12'h333;
			{8'd140, 8'd96}: color_data = 12'h333;
			{8'd140, 8'd97}: color_data = 12'h333;
			{8'd140, 8'd98}: color_data = 12'h333;
			{8'd140, 8'd99}: color_data = 12'h333;
			{8'd140, 8'd100}: color_data = 12'h333;
			{8'd140, 8'd101}: color_data = 12'h333;
			{8'd140, 8'd102}: color_data = 12'h333;
			{8'd140, 8'd103}: color_data = 12'h333;
			{8'd140, 8'd104}: color_data = 12'h333;
			{8'd140, 8'd105}: color_data = 12'h333;
			{8'd140, 8'd106}: color_data = 12'h333;
			{8'd140, 8'd107}: color_data = 12'h222;
			{8'd140, 8'd108}: color_data = 12'h222;
			{8'd140, 8'd109}: color_data = 12'h222;
			{8'd140, 8'd110}: color_data = 12'h222;
			{8'd140, 8'd111}: color_data = 12'h222;
			{8'd140, 8'd112}: color_data = 12'h222;
			{8'd140, 8'd113}: color_data = 12'h222;
			{8'd140, 8'd114}: color_data = 12'h222;
			{8'd140, 8'd115}: color_data = 12'h222;
			{8'd140, 8'd116}: color_data = 12'h222;
			{8'd140, 8'd117}: color_data = 12'h222;
			{8'd140, 8'd118}: color_data = 12'h222;
			{8'd140, 8'd119}: color_data = 12'h222;
			{8'd140, 8'd120}: color_data = 12'h222;
			{8'd140, 8'd121}: color_data = 12'h111;
			{8'd140, 8'd122}: color_data = 12'h111;
			{8'd140, 8'd123}: color_data = 12'h111;
			{8'd140, 8'd124}: color_data = 12'h222;
			{8'd140, 8'd125}: color_data = 12'haaa;
			{8'd140, 8'd126}: color_data = 12'hfff;
			{8'd140, 8'd127}: color_data = 12'hfff;
			{8'd140, 8'd128}: color_data = 12'hfff;
			{8'd140, 8'd129}: color_data = 12'hfff;
			{8'd140, 8'd130}: color_data = 12'hfff;
			{8'd140, 8'd131}: color_data = 12'hfff;
			{8'd140, 8'd132}: color_data = 12'hfff;
			{8'd140, 8'd133}: color_data = 12'hfff;
			{8'd140, 8'd134}: color_data = 12'hfff;
			{8'd140, 8'd135}: color_data = 12'hfff;
			{8'd140, 8'd136}: color_data = 12'hfff;
			{8'd140, 8'd137}: color_data = 12'heee;
			{8'd140, 8'd138}: color_data = 12'h888;
			{8'd140, 8'd139}: color_data = 12'h555;
			{8'd141, 8'd32}: color_data = 12'hb11;
			{8'd141, 8'd33}: color_data = 12'hd11;
			{8'd141, 8'd34}: color_data = 12'hd21;
			{8'd141, 8'd35}: color_data = 12'hd21;
			{8'd141, 8'd36}: color_data = 12'hd31;
			{8'd141, 8'd37}: color_data = 12'hb31;
			{8'd141, 8'd38}: color_data = 12'h920;
			{8'd141, 8'd44}: color_data = 12'h730;
			{8'd141, 8'd45}: color_data = 12'hb50;
			{8'd141, 8'd46}: color_data = 12'hd70;
			{8'd141, 8'd47}: color_data = 12'he80;
			{8'd141, 8'd48}: color_data = 12'he80;
			{8'd141, 8'd49}: color_data = 12'he80;
			{8'd141, 8'd50}: color_data = 12'he90;
			{8'd141, 8'd51}: color_data = 12'he90;
			{8'd141, 8'd52}: color_data = 12'hd80;
			{8'd141, 8'd53}: color_data = 12'ha70;
			{8'd141, 8'd60}: color_data = 12'h999;
			{8'd141, 8'd61}: color_data = 12'h666;
			{8'd141, 8'd62}: color_data = 12'h555;
			{8'd141, 8'd63}: color_data = 12'h666;
			{8'd141, 8'd64}: color_data = 12'h666;
			{8'd141, 8'd65}: color_data = 12'h666;
			{8'd141, 8'd66}: color_data = 12'h666;
			{8'd141, 8'd67}: color_data = 12'h666;
			{8'd141, 8'd68}: color_data = 12'h555;
			{8'd141, 8'd69}: color_data = 12'h555;
			{8'd141, 8'd70}: color_data = 12'h555;
			{8'd141, 8'd71}: color_data = 12'h555;
			{8'd141, 8'd72}: color_data = 12'h555;
			{8'd141, 8'd73}: color_data = 12'h555;
			{8'd141, 8'd74}: color_data = 12'h555;
			{8'd141, 8'd75}: color_data = 12'h555;
			{8'd141, 8'd76}: color_data = 12'h555;
			{8'd141, 8'd77}: color_data = 12'h555;
			{8'd141, 8'd78}: color_data = 12'h555;
			{8'd141, 8'd79}: color_data = 12'h555;
			{8'd141, 8'd80}: color_data = 12'h444;
			{8'd141, 8'd81}: color_data = 12'h444;
			{8'd141, 8'd82}: color_data = 12'h444;
			{8'd141, 8'd83}: color_data = 12'h444;
			{8'd141, 8'd84}: color_data = 12'h444;
			{8'd141, 8'd85}: color_data = 12'h444;
			{8'd141, 8'd86}: color_data = 12'h444;
			{8'd141, 8'd87}: color_data = 12'h444;
			{8'd141, 8'd88}: color_data = 12'h444;
			{8'd141, 8'd89}: color_data = 12'h444;
			{8'd141, 8'd90}: color_data = 12'h444;
			{8'd141, 8'd91}: color_data = 12'h444;
			{8'd141, 8'd92}: color_data = 12'h444;
			{8'd141, 8'd93}: color_data = 12'h444;
			{8'd141, 8'd94}: color_data = 12'h333;
			{8'd141, 8'd95}: color_data = 12'h333;
			{8'd141, 8'd96}: color_data = 12'h333;
			{8'd141, 8'd97}: color_data = 12'h333;
			{8'd141, 8'd98}: color_data = 12'h333;
			{8'd141, 8'd99}: color_data = 12'h333;
			{8'd141, 8'd100}: color_data = 12'h333;
			{8'd141, 8'd101}: color_data = 12'h333;
			{8'd141, 8'd102}: color_data = 12'h333;
			{8'd141, 8'd103}: color_data = 12'h333;
			{8'd141, 8'd104}: color_data = 12'h333;
			{8'd141, 8'd105}: color_data = 12'h333;
			{8'd141, 8'd106}: color_data = 12'h333;
			{8'd141, 8'd107}: color_data = 12'h222;
			{8'd141, 8'd108}: color_data = 12'h222;
			{8'd141, 8'd109}: color_data = 12'h222;
			{8'd141, 8'd110}: color_data = 12'h222;
			{8'd141, 8'd111}: color_data = 12'h222;
			{8'd141, 8'd112}: color_data = 12'h222;
			{8'd141, 8'd113}: color_data = 12'h222;
			{8'd141, 8'd114}: color_data = 12'h222;
			{8'd141, 8'd115}: color_data = 12'h222;
			{8'd141, 8'd116}: color_data = 12'h222;
			{8'd141, 8'd117}: color_data = 12'h222;
			{8'd141, 8'd118}: color_data = 12'h222;
			{8'd141, 8'd119}: color_data = 12'h222;
			{8'd141, 8'd120}: color_data = 12'h222;
			{8'd141, 8'd121}: color_data = 12'h111;
			{8'd141, 8'd122}: color_data = 12'h111;
			{8'd141, 8'd123}: color_data = 12'h111;
			{8'd141, 8'd124}: color_data = 12'h111;
			{8'd141, 8'd125}: color_data = 12'h777;
			{8'd141, 8'd126}: color_data = 12'heee;
			{8'd141, 8'd127}: color_data = 12'hfff;
			{8'd141, 8'd128}: color_data = 12'hfff;
			{8'd141, 8'd129}: color_data = 12'hfff;
			{8'd141, 8'd130}: color_data = 12'hfff;
			{8'd141, 8'd131}: color_data = 12'hfff;
			{8'd141, 8'd132}: color_data = 12'hfff;
			{8'd141, 8'd133}: color_data = 12'hfff;
			{8'd141, 8'd134}: color_data = 12'hfff;
			{8'd141, 8'd135}: color_data = 12'hfff;
			{8'd141, 8'd136}: color_data = 12'hfff;
			{8'd141, 8'd137}: color_data = 12'hddd;
			{8'd141, 8'd138}: color_data = 12'h777;
			{8'd141, 8'd139}: color_data = 12'h444;
			{8'd142, 8'd32}: color_data = 12'ha11;
			{8'd142, 8'd33}: color_data = 12'hc11;
			{8'd142, 8'd34}: color_data = 12'hd21;
			{8'd142, 8'd35}: color_data = 12'hd21;
			{8'd142, 8'd36}: color_data = 12'hd31;
			{8'd142, 8'd37}: color_data = 12'hd31;
			{8'd142, 8'd38}: color_data = 12'hb31;
			{8'd142, 8'd39}: color_data = 12'ha30;
			{8'd142, 8'd40}: color_data = 12'hc41;
			{8'd142, 8'd41}: color_data = 12'hc41;
			{8'd142, 8'd42}: color_data = 12'hc50;
			{8'd142, 8'd43}: color_data = 12'hc51;
			{8'd142, 8'd44}: color_data = 12'hb50;
			{8'd142, 8'd45}: color_data = 12'hc61;
			{8'd142, 8'd46}: color_data = 12'he71;
			{8'd142, 8'd47}: color_data = 12'he80;
			{8'd142, 8'd48}: color_data = 12'he80;
			{8'd142, 8'd49}: color_data = 12'he80;
			{8'd142, 8'd50}: color_data = 12'he90;
			{8'd142, 8'd51}: color_data = 12'he90;
			{8'd142, 8'd52}: color_data = 12'hb70;
			{8'd142, 8'd53}: color_data = 12'h950;
			{8'd142, 8'd66}: color_data = 12'h555;
			{8'd142, 8'd67}: color_data = 12'h555;
			{8'd142, 8'd68}: color_data = 12'h555;
			{8'd142, 8'd69}: color_data = 12'h555;
			{8'd142, 8'd70}: color_data = 12'h555;
			{8'd142, 8'd71}: color_data = 12'h555;
			{8'd142, 8'd72}: color_data = 12'h555;
			{8'd142, 8'd73}: color_data = 12'h555;
			{8'd142, 8'd74}: color_data = 12'h555;
			{8'd142, 8'd75}: color_data = 12'h555;
			{8'd142, 8'd76}: color_data = 12'h555;
			{8'd142, 8'd77}: color_data = 12'h555;
			{8'd142, 8'd78}: color_data = 12'h555;
			{8'd142, 8'd79}: color_data = 12'h555;
			{8'd142, 8'd80}: color_data = 12'h444;
			{8'd142, 8'd81}: color_data = 12'h444;
			{8'd142, 8'd82}: color_data = 12'h444;
			{8'd142, 8'd83}: color_data = 12'h444;
			{8'd142, 8'd84}: color_data = 12'h444;
			{8'd142, 8'd85}: color_data = 12'h444;
			{8'd142, 8'd86}: color_data = 12'h444;
			{8'd142, 8'd87}: color_data = 12'h444;
			{8'd142, 8'd88}: color_data = 12'h444;
			{8'd142, 8'd89}: color_data = 12'h444;
			{8'd142, 8'd90}: color_data = 12'h444;
			{8'd142, 8'd91}: color_data = 12'h444;
			{8'd142, 8'd92}: color_data = 12'h444;
			{8'd142, 8'd93}: color_data = 12'h444;
			{8'd142, 8'd94}: color_data = 12'h333;
			{8'd142, 8'd95}: color_data = 12'h333;
			{8'd142, 8'd96}: color_data = 12'h333;
			{8'd142, 8'd97}: color_data = 12'h333;
			{8'd142, 8'd98}: color_data = 12'h333;
			{8'd142, 8'd99}: color_data = 12'h333;
			{8'd142, 8'd100}: color_data = 12'h333;
			{8'd142, 8'd101}: color_data = 12'h333;
			{8'd142, 8'd102}: color_data = 12'h333;
			{8'd142, 8'd103}: color_data = 12'h333;
			{8'd142, 8'd104}: color_data = 12'h333;
			{8'd142, 8'd105}: color_data = 12'h333;
			{8'd142, 8'd106}: color_data = 12'h333;
			{8'd142, 8'd107}: color_data = 12'h222;
			{8'd142, 8'd108}: color_data = 12'h222;
			{8'd142, 8'd109}: color_data = 12'h222;
			{8'd142, 8'd110}: color_data = 12'h222;
			{8'd142, 8'd111}: color_data = 12'h222;
			{8'd142, 8'd112}: color_data = 12'h222;
			{8'd142, 8'd113}: color_data = 12'h222;
			{8'd142, 8'd114}: color_data = 12'h222;
			{8'd142, 8'd115}: color_data = 12'h222;
			{8'd142, 8'd116}: color_data = 12'h222;
			{8'd142, 8'd117}: color_data = 12'h222;
			{8'd142, 8'd118}: color_data = 12'h222;
			{8'd142, 8'd119}: color_data = 12'h222;
			{8'd142, 8'd120}: color_data = 12'h111;
			{8'd142, 8'd121}: color_data = 12'h111;
			{8'd142, 8'd122}: color_data = 12'h111;
			{8'd142, 8'd123}: color_data = 12'h111;
			{8'd142, 8'd124}: color_data = 12'h111;
			{8'd142, 8'd125}: color_data = 12'h555;
			{8'd142, 8'd126}: color_data = 12'hddd;
			{8'd142, 8'd127}: color_data = 12'hfff;
			{8'd142, 8'd128}: color_data = 12'hfff;
			{8'd142, 8'd129}: color_data = 12'hfff;
			{8'd142, 8'd130}: color_data = 12'hfff;
			{8'd142, 8'd131}: color_data = 12'hfff;
			{8'd142, 8'd132}: color_data = 12'hfff;
			{8'd142, 8'd133}: color_data = 12'hfff;
			{8'd142, 8'd134}: color_data = 12'hfff;
			{8'd142, 8'd135}: color_data = 12'hfff;
			{8'd142, 8'd136}: color_data = 12'hfff;
			{8'd142, 8'd137}: color_data = 12'hbbb;
			{8'd142, 8'd138}: color_data = 12'h777;
			{8'd143, 8'd32}: color_data = 12'h700;
			{8'd143, 8'd33}: color_data = 12'hb11;
			{8'd143, 8'd34}: color_data = 12'hd21;
			{8'd143, 8'd35}: color_data = 12'hd21;
			{8'd143, 8'd36}: color_data = 12'hd31;
			{8'd143, 8'd37}: color_data = 12'he41;
			{8'd143, 8'd38}: color_data = 12'hd41;
			{8'd143, 8'd39}: color_data = 12'hc41;
			{8'd143, 8'd40}: color_data = 12'hc41;
			{8'd143, 8'd41}: color_data = 12'hc51;
			{8'd143, 8'd42}: color_data = 12'hc51;
			{8'd143, 8'd43}: color_data = 12'hc51;
			{8'd143, 8'd44}: color_data = 12'hd61;
			{8'd143, 8'd45}: color_data = 12'he71;
			{8'd143, 8'd46}: color_data = 12'he71;
			{8'd143, 8'd47}: color_data = 12'he80;
			{8'd143, 8'd48}: color_data = 12'he80;
			{8'd143, 8'd49}: color_data = 12'he80;
			{8'd143, 8'd50}: color_data = 12'he80;
			{8'd143, 8'd51}: color_data = 12'hc80;
			{8'd143, 8'd52}: color_data = 12'h960;
			{8'd143, 8'd70}: color_data = 12'h000;
			{8'd143, 8'd71}: color_data = 12'h333;
			{8'd143, 8'd72}: color_data = 12'h555;
			{8'd143, 8'd73}: color_data = 12'h555;
			{8'd143, 8'd74}: color_data = 12'h555;
			{8'd143, 8'd75}: color_data = 12'h555;
			{8'd143, 8'd76}: color_data = 12'h555;
			{8'd143, 8'd77}: color_data = 12'h555;
			{8'd143, 8'd78}: color_data = 12'h555;
			{8'd143, 8'd79}: color_data = 12'h444;
			{8'd143, 8'd80}: color_data = 12'h444;
			{8'd143, 8'd81}: color_data = 12'h555;
			{8'd143, 8'd82}: color_data = 12'h444;
			{8'd143, 8'd83}: color_data = 12'h444;
			{8'd143, 8'd84}: color_data = 12'h444;
			{8'd143, 8'd85}: color_data = 12'h444;
			{8'd143, 8'd86}: color_data = 12'h444;
			{8'd143, 8'd87}: color_data = 12'h444;
			{8'd143, 8'd88}: color_data = 12'h444;
			{8'd143, 8'd89}: color_data = 12'h444;
			{8'd143, 8'd90}: color_data = 12'h444;
			{8'd143, 8'd91}: color_data = 12'h444;
			{8'd143, 8'd92}: color_data = 12'h444;
			{8'd143, 8'd93}: color_data = 12'h333;
			{8'd143, 8'd94}: color_data = 12'h333;
			{8'd143, 8'd95}: color_data = 12'h333;
			{8'd143, 8'd96}: color_data = 12'h333;
			{8'd143, 8'd97}: color_data = 12'h333;
			{8'd143, 8'd98}: color_data = 12'h333;
			{8'd143, 8'd99}: color_data = 12'h333;
			{8'd143, 8'd100}: color_data = 12'h333;
			{8'd143, 8'd101}: color_data = 12'h333;
			{8'd143, 8'd102}: color_data = 12'h333;
			{8'd143, 8'd103}: color_data = 12'h333;
			{8'd143, 8'd104}: color_data = 12'h333;
			{8'd143, 8'd105}: color_data = 12'h333;
			{8'd143, 8'd106}: color_data = 12'h222;
			{8'd143, 8'd107}: color_data = 12'h222;
			{8'd143, 8'd108}: color_data = 12'h222;
			{8'd143, 8'd109}: color_data = 12'h222;
			{8'd143, 8'd110}: color_data = 12'h222;
			{8'd143, 8'd111}: color_data = 12'h222;
			{8'd143, 8'd112}: color_data = 12'h222;
			{8'd143, 8'd113}: color_data = 12'h222;
			{8'd143, 8'd114}: color_data = 12'h222;
			{8'd143, 8'd115}: color_data = 12'h222;
			{8'd143, 8'd116}: color_data = 12'h222;
			{8'd143, 8'd117}: color_data = 12'h222;
			{8'd143, 8'd118}: color_data = 12'h222;
			{8'd143, 8'd119}: color_data = 12'h222;
			{8'd143, 8'd120}: color_data = 12'h111;
			{8'd143, 8'd121}: color_data = 12'h111;
			{8'd143, 8'd122}: color_data = 12'h111;
			{8'd143, 8'd123}: color_data = 12'h111;
			{8'd143, 8'd124}: color_data = 12'h111;
			{8'd143, 8'd125}: color_data = 12'h333;
			{8'd143, 8'd126}: color_data = 12'haaa;
			{8'd143, 8'd127}: color_data = 12'hfff;
			{8'd143, 8'd128}: color_data = 12'hfff;
			{8'd143, 8'd129}: color_data = 12'hfff;
			{8'd143, 8'd130}: color_data = 12'hfff;
			{8'd143, 8'd131}: color_data = 12'hfff;
			{8'd143, 8'd132}: color_data = 12'hfff;
			{8'd143, 8'd133}: color_data = 12'hfff;
			{8'd143, 8'd134}: color_data = 12'hfff;
			{8'd143, 8'd135}: color_data = 12'hfff;
			{8'd143, 8'd136}: color_data = 12'heee;
			{8'd143, 8'd137}: color_data = 12'h999;
			{8'd143, 8'd138}: color_data = 12'h666;
			{8'd144, 8'd33}: color_data = 12'ha11;
			{8'd144, 8'd34}: color_data = 12'hb21;
			{8'd144, 8'd35}: color_data = 12'hd21;
			{8'd144, 8'd36}: color_data = 12'he31;
			{8'd144, 8'd37}: color_data = 12'hd41;
			{8'd144, 8'd38}: color_data = 12'he41;
			{8'd144, 8'd39}: color_data = 12'he51;
			{8'd144, 8'd40}: color_data = 12'he51;
			{8'd144, 8'd41}: color_data = 12'he51;
			{8'd144, 8'd42}: color_data = 12'he61;
			{8'd144, 8'd43}: color_data = 12'he61;
			{8'd144, 8'd44}: color_data = 12'he71;
			{8'd144, 8'd45}: color_data = 12'he71;
			{8'd144, 8'd46}: color_data = 12'he71;
			{8'd144, 8'd47}: color_data = 12'he80;
			{8'd144, 8'd48}: color_data = 12'he80;
			{8'd144, 8'd49}: color_data = 12'he80;
			{8'd144, 8'd50}: color_data = 12'hc70;
			{8'd144, 8'd51}: color_data = 12'ha60;
			{8'd144, 8'd76}: color_data = 12'h555;
			{8'd144, 8'd77}: color_data = 12'h555;
			{8'd144, 8'd78}: color_data = 12'h555;
			{8'd144, 8'd79}: color_data = 12'h444;
			{8'd144, 8'd80}: color_data = 12'h444;
			{8'd144, 8'd81}: color_data = 12'h444;
			{8'd144, 8'd82}: color_data = 12'h444;
			{8'd144, 8'd83}: color_data = 12'h444;
			{8'd144, 8'd84}: color_data = 12'h444;
			{8'd144, 8'd85}: color_data = 12'h444;
			{8'd144, 8'd86}: color_data = 12'h444;
			{8'd144, 8'd87}: color_data = 12'h444;
			{8'd144, 8'd88}: color_data = 12'h444;
			{8'd144, 8'd89}: color_data = 12'h444;
			{8'd144, 8'd90}: color_data = 12'h444;
			{8'd144, 8'd91}: color_data = 12'h444;
			{8'd144, 8'd92}: color_data = 12'h333;
			{8'd144, 8'd93}: color_data = 12'h333;
			{8'd144, 8'd94}: color_data = 12'h333;
			{8'd144, 8'd95}: color_data = 12'h333;
			{8'd144, 8'd96}: color_data = 12'h333;
			{8'd144, 8'd97}: color_data = 12'h333;
			{8'd144, 8'd98}: color_data = 12'h333;
			{8'd144, 8'd99}: color_data = 12'h333;
			{8'd144, 8'd100}: color_data = 12'h333;
			{8'd144, 8'd101}: color_data = 12'h333;
			{8'd144, 8'd102}: color_data = 12'h333;
			{8'd144, 8'd103}: color_data = 12'h333;
			{8'd144, 8'd104}: color_data = 12'h333;
			{8'd144, 8'd105}: color_data = 12'h222;
			{8'd144, 8'd106}: color_data = 12'h222;
			{8'd144, 8'd107}: color_data = 12'h222;
			{8'd144, 8'd108}: color_data = 12'h222;
			{8'd144, 8'd109}: color_data = 12'h222;
			{8'd144, 8'd110}: color_data = 12'h222;
			{8'd144, 8'd111}: color_data = 12'h222;
			{8'd144, 8'd112}: color_data = 12'h222;
			{8'd144, 8'd113}: color_data = 12'h222;
			{8'd144, 8'd114}: color_data = 12'h222;
			{8'd144, 8'd115}: color_data = 12'h222;
			{8'd144, 8'd116}: color_data = 12'h222;
			{8'd144, 8'd117}: color_data = 12'h222;
			{8'd144, 8'd118}: color_data = 12'h222;
			{8'd144, 8'd119}: color_data = 12'h111;
			{8'd144, 8'd120}: color_data = 12'h111;
			{8'd144, 8'd121}: color_data = 12'h111;
			{8'd144, 8'd122}: color_data = 12'h111;
			{8'd144, 8'd123}: color_data = 12'h111;
			{8'd144, 8'd124}: color_data = 12'h111;
			{8'd144, 8'd125}: color_data = 12'h222;
			{8'd144, 8'd126}: color_data = 12'h777;
			{8'd144, 8'd127}: color_data = 12'heee;
			{8'd144, 8'd128}: color_data = 12'hfff;
			{8'd144, 8'd129}: color_data = 12'hfff;
			{8'd144, 8'd130}: color_data = 12'hfff;
			{8'd144, 8'd131}: color_data = 12'hfff;
			{8'd144, 8'd132}: color_data = 12'hfff;
			{8'd144, 8'd133}: color_data = 12'hfff;
			{8'd144, 8'd134}: color_data = 12'hfff;
			{8'd144, 8'd135}: color_data = 12'hfff;
			{8'd144, 8'd136}: color_data = 12'hddd;
			{8'd144, 8'd137}: color_data = 12'h888;
			{8'd144, 8'd138}: color_data = 12'h111;
			{8'd145, 8'd34}: color_data = 12'h910;
			{8'd145, 8'd35}: color_data = 12'hb21;
			{8'd145, 8'd36}: color_data = 12'hc31;
			{8'd145, 8'd37}: color_data = 12'he41;
			{8'd145, 8'd38}: color_data = 12'he41;
			{8'd145, 8'd39}: color_data = 12'he51;
			{8'd145, 8'd40}: color_data = 12'he51;
			{8'd145, 8'd41}: color_data = 12'he51;
			{8'd145, 8'd42}: color_data = 12'he61;
			{8'd145, 8'd43}: color_data = 12'he61;
			{8'd145, 8'd44}: color_data = 12'he71;
			{8'd145, 8'd45}: color_data = 12'he71;
			{8'd145, 8'd46}: color_data = 12'he71;
			{8'd145, 8'd47}: color_data = 12'he80;
			{8'd145, 8'd48}: color_data = 12'he80;
			{8'd145, 8'd49}: color_data = 12'hc70;
			{8'd145, 8'd50}: color_data = 12'ha60;
			{8'd145, 8'd82}: color_data = 12'h444;
			{8'd145, 8'd83}: color_data = 12'h444;
			{8'd145, 8'd84}: color_data = 12'h444;
			{8'd145, 8'd85}: color_data = 12'h444;
			{8'd145, 8'd86}: color_data = 12'h444;
			{8'd145, 8'd87}: color_data = 12'h444;
			{8'd145, 8'd88}: color_data = 12'h444;
			{8'd145, 8'd89}: color_data = 12'h444;
			{8'd145, 8'd90}: color_data = 12'h444;
			{8'd145, 8'd91}: color_data = 12'h444;
			{8'd145, 8'd92}: color_data = 12'h444;
			{8'd145, 8'd93}: color_data = 12'h444;
			{8'd145, 8'd94}: color_data = 12'h333;
			{8'd145, 8'd95}: color_data = 12'h333;
			{8'd145, 8'd96}: color_data = 12'h333;
			{8'd145, 8'd97}: color_data = 12'h333;
			{8'd145, 8'd98}: color_data = 12'h333;
			{8'd145, 8'd99}: color_data = 12'h333;
			{8'd145, 8'd100}: color_data = 12'h333;
			{8'd145, 8'd101}: color_data = 12'h333;
			{8'd145, 8'd102}: color_data = 12'h333;
			{8'd145, 8'd103}: color_data = 12'h333;
			{8'd145, 8'd104}: color_data = 12'h333;
			{8'd145, 8'd105}: color_data = 12'h333;
			{8'd145, 8'd106}: color_data = 12'h222;
			{8'd145, 8'd107}: color_data = 12'h222;
			{8'd145, 8'd108}: color_data = 12'h222;
			{8'd145, 8'd109}: color_data = 12'h222;
			{8'd145, 8'd110}: color_data = 12'h222;
			{8'd145, 8'd111}: color_data = 12'h222;
			{8'd145, 8'd112}: color_data = 12'h222;
			{8'd145, 8'd113}: color_data = 12'h222;
			{8'd145, 8'd114}: color_data = 12'h222;
			{8'd145, 8'd115}: color_data = 12'h222;
			{8'd145, 8'd116}: color_data = 12'h222;
			{8'd145, 8'd117}: color_data = 12'h222;
			{8'd145, 8'd118}: color_data = 12'h222;
			{8'd145, 8'd119}: color_data = 12'h111;
			{8'd145, 8'd120}: color_data = 12'h111;
			{8'd145, 8'd121}: color_data = 12'h111;
			{8'd145, 8'd122}: color_data = 12'h111;
			{8'd145, 8'd123}: color_data = 12'h111;
			{8'd145, 8'd124}: color_data = 12'h111;
			{8'd145, 8'd125}: color_data = 12'h111;
			{8'd145, 8'd126}: color_data = 12'h444;
			{8'd145, 8'd127}: color_data = 12'hccc;
			{8'd145, 8'd128}: color_data = 12'hfff;
			{8'd145, 8'd129}: color_data = 12'hfff;
			{8'd145, 8'd130}: color_data = 12'hfff;
			{8'd145, 8'd131}: color_data = 12'hfff;
			{8'd145, 8'd132}: color_data = 12'hfff;
			{8'd145, 8'd133}: color_data = 12'hfff;
			{8'd145, 8'd134}: color_data = 12'hfff;
			{8'd145, 8'd135}: color_data = 12'heee;
			{8'd145, 8'd136}: color_data = 12'haaa;
			{8'd145, 8'd137}: color_data = 12'h666;
			{8'd146, 8'd35}: color_data = 12'h721;
			{8'd146, 8'd36}: color_data = 12'ha20;
			{8'd146, 8'd37}: color_data = 12'hd31;
			{8'd146, 8'd38}: color_data = 12'he41;
			{8'd146, 8'd39}: color_data = 12'he51;
			{8'd146, 8'd40}: color_data = 12'he51;
			{8'd146, 8'd41}: color_data = 12'he61;
			{8'd146, 8'd42}: color_data = 12'he61;
			{8'd146, 8'd43}: color_data = 12'he61;
			{8'd146, 8'd44}: color_data = 12'he71;
			{8'd146, 8'd45}: color_data = 12'he71;
			{8'd146, 8'd46}: color_data = 12'he71;
			{8'd146, 8'd47}: color_data = 12'he80;
			{8'd146, 8'd48}: color_data = 12'hc70;
			{8'd146, 8'd49}: color_data = 12'hb60;
			{8'd146, 8'd86}: color_data = 12'h000;
			{8'd146, 8'd87}: color_data = 12'h444;
			{8'd146, 8'd88}: color_data = 12'h444;
			{8'd146, 8'd89}: color_data = 12'h444;
			{8'd146, 8'd90}: color_data = 12'h333;
			{8'd146, 8'd91}: color_data = 12'h333;
			{8'd146, 8'd92}: color_data = 12'h333;
			{8'd146, 8'd93}: color_data = 12'h333;
			{8'd146, 8'd94}: color_data = 12'h333;
			{8'd146, 8'd95}: color_data = 12'h333;
			{8'd146, 8'd96}: color_data = 12'h333;
			{8'd146, 8'd97}: color_data = 12'h333;
			{8'd146, 8'd98}: color_data = 12'h333;
			{8'd146, 8'd99}: color_data = 12'h333;
			{8'd146, 8'd100}: color_data = 12'h333;
			{8'd146, 8'd101}: color_data = 12'h333;
			{8'd146, 8'd102}: color_data = 12'h333;
			{8'd146, 8'd103}: color_data = 12'h333;
			{8'd146, 8'd104}: color_data = 12'h222;
			{8'd146, 8'd105}: color_data = 12'h222;
			{8'd146, 8'd106}: color_data = 12'h222;
			{8'd146, 8'd107}: color_data = 12'h222;
			{8'd146, 8'd108}: color_data = 12'h222;
			{8'd146, 8'd109}: color_data = 12'h222;
			{8'd146, 8'd110}: color_data = 12'h222;
			{8'd146, 8'd111}: color_data = 12'h222;
			{8'd146, 8'd112}: color_data = 12'h222;
			{8'd146, 8'd113}: color_data = 12'h222;
			{8'd146, 8'd114}: color_data = 12'h222;
			{8'd146, 8'd115}: color_data = 12'h222;
			{8'd146, 8'd116}: color_data = 12'h222;
			{8'd146, 8'd117}: color_data = 12'h222;
			{8'd146, 8'd118}: color_data = 12'h111;
			{8'd146, 8'd119}: color_data = 12'h111;
			{8'd146, 8'd120}: color_data = 12'h111;
			{8'd146, 8'd121}: color_data = 12'h111;
			{8'd146, 8'd122}: color_data = 12'h111;
			{8'd146, 8'd123}: color_data = 12'h111;
			{8'd146, 8'd124}: color_data = 12'h111;
			{8'd146, 8'd125}: color_data = 12'h111;
			{8'd146, 8'd126}: color_data = 12'h222;
			{8'd146, 8'd127}: color_data = 12'h999;
			{8'd146, 8'd128}: color_data = 12'heee;
			{8'd146, 8'd129}: color_data = 12'hfff;
			{8'd146, 8'd130}: color_data = 12'hfff;
			{8'd146, 8'd131}: color_data = 12'hfff;
			{8'd146, 8'd132}: color_data = 12'hfff;
			{8'd146, 8'd133}: color_data = 12'hfff;
			{8'd146, 8'd134}: color_data = 12'hfff;
			{8'd146, 8'd135}: color_data = 12'hddd;
			{8'd146, 8'd136}: color_data = 12'h888;
			{8'd146, 8'd137}: color_data = 12'h555;
			{8'd147, 8'd36}: color_data = 12'h821;
			{8'd147, 8'd37}: color_data = 12'ha30;
			{8'd147, 8'd38}: color_data = 12'hc41;
			{8'd147, 8'd39}: color_data = 12'hd41;
			{8'd147, 8'd40}: color_data = 12'he51;
			{8'd147, 8'd41}: color_data = 12'he51;
			{8'd147, 8'd42}: color_data = 12'he61;
			{8'd147, 8'd43}: color_data = 12'he61;
			{8'd147, 8'd44}: color_data = 12'he61;
			{8'd147, 8'd45}: color_data = 12'hd71;
			{8'd147, 8'd46}: color_data = 12'hd71;
			{8'd147, 8'd47}: color_data = 12'hd70;
			{8'd147, 8'd48}: color_data = 12'hc70;
			{8'd147, 8'd91}: color_data = 12'h333;
			{8'd147, 8'd92}: color_data = 12'h555;
			{8'd147, 8'd93}: color_data = 12'h333;
			{8'd147, 8'd94}: color_data = 12'h333;
			{8'd147, 8'd95}: color_data = 12'h333;
			{8'd147, 8'd96}: color_data = 12'h333;
			{8'd147, 8'd97}: color_data = 12'h333;
			{8'd147, 8'd98}: color_data = 12'h333;
			{8'd147, 8'd99}: color_data = 12'h333;
			{8'd147, 8'd100}: color_data = 12'h333;
			{8'd147, 8'd101}: color_data = 12'h333;
			{8'd147, 8'd102}: color_data = 12'h333;
			{8'd147, 8'd103}: color_data = 12'h333;
			{8'd147, 8'd104}: color_data = 12'h333;
			{8'd147, 8'd105}: color_data = 12'h333;
			{8'd147, 8'd106}: color_data = 12'h222;
			{8'd147, 8'd107}: color_data = 12'h222;
			{8'd147, 8'd108}: color_data = 12'h222;
			{8'd147, 8'd109}: color_data = 12'h222;
			{8'd147, 8'd110}: color_data = 12'h222;
			{8'd147, 8'd111}: color_data = 12'h222;
			{8'd147, 8'd112}: color_data = 12'h222;
			{8'd147, 8'd113}: color_data = 12'h222;
			{8'd147, 8'd114}: color_data = 12'h222;
			{8'd147, 8'd115}: color_data = 12'h222;
			{8'd147, 8'd116}: color_data = 12'h222;
			{8'd147, 8'd117}: color_data = 12'h222;
			{8'd147, 8'd118}: color_data = 12'h111;
			{8'd147, 8'd119}: color_data = 12'h111;
			{8'd147, 8'd120}: color_data = 12'h111;
			{8'd147, 8'd121}: color_data = 12'h111;
			{8'd147, 8'd122}: color_data = 12'h111;
			{8'd147, 8'd123}: color_data = 12'h111;
			{8'd147, 8'd124}: color_data = 12'h111;
			{8'd147, 8'd125}: color_data = 12'h111;
			{8'd147, 8'd126}: color_data = 12'h111;
			{8'd147, 8'd127}: color_data = 12'h555;
			{8'd147, 8'd128}: color_data = 12'hccc;
			{8'd147, 8'd129}: color_data = 12'heee;
			{8'd147, 8'd130}: color_data = 12'hfff;
			{8'd147, 8'd131}: color_data = 12'hfff;
			{8'd147, 8'd132}: color_data = 12'hfff;
			{8'd147, 8'd133}: color_data = 12'hfff;
			{8'd147, 8'd134}: color_data = 12'heee;
			{8'd147, 8'd135}: color_data = 12'haaa;
			{8'd147, 8'd136}: color_data = 12'h666;
			{8'd147, 8'd137}: color_data = 12'h555;
			{8'd148, 8'd37}: color_data = 12'h720;
			{8'd148, 8'd38}: color_data = 12'h920;
			{8'd148, 8'd39}: color_data = 12'hc41;
			{8'd148, 8'd40}: color_data = 12'hd51;
			{8'd148, 8'd41}: color_data = 12'hd61;
			{8'd148, 8'd42}: color_data = 12'hd61;
			{8'd148, 8'd43}: color_data = 12'hd61;
			{8'd148, 8'd44}: color_data = 12'hd61;
			{8'd148, 8'd45}: color_data = 12'hd71;
			{8'd148, 8'd46}: color_data = 12'hd61;
			{8'd148, 8'd47}: color_data = 12'he61;
			{8'd148, 8'd97}: color_data = 12'h333;
			{8'd148, 8'd98}: color_data = 12'h333;
			{8'd148, 8'd99}: color_data = 12'h333;
			{8'd148, 8'd100}: color_data = 12'h333;
			{8'd148, 8'd101}: color_data = 12'h333;
			{8'd148, 8'd102}: color_data = 12'h333;
			{8'd148, 8'd103}: color_data = 12'h222;
			{8'd148, 8'd104}: color_data = 12'h222;
			{8'd148, 8'd105}: color_data = 12'h222;
			{8'd148, 8'd106}: color_data = 12'h222;
			{8'd148, 8'd107}: color_data = 12'h222;
			{8'd148, 8'd108}: color_data = 12'h222;
			{8'd148, 8'd109}: color_data = 12'h222;
			{8'd148, 8'd110}: color_data = 12'h222;
			{8'd148, 8'd111}: color_data = 12'h222;
			{8'd148, 8'd112}: color_data = 12'h222;
			{8'd148, 8'd113}: color_data = 12'h222;
			{8'd148, 8'd114}: color_data = 12'h222;
			{8'd148, 8'd115}: color_data = 12'h222;
			{8'd148, 8'd116}: color_data = 12'h222;
			{8'd148, 8'd117}: color_data = 12'h222;
			{8'd148, 8'd118}: color_data = 12'h111;
			{8'd148, 8'd119}: color_data = 12'h111;
			{8'd148, 8'd120}: color_data = 12'h111;
			{8'd148, 8'd121}: color_data = 12'h111;
			{8'd148, 8'd122}: color_data = 12'h111;
			{8'd148, 8'd123}: color_data = 12'h111;
			{8'd148, 8'd124}: color_data = 12'h111;
			{8'd148, 8'd125}: color_data = 12'h111;
			{8'd148, 8'd126}: color_data = 12'h111;
			{8'd148, 8'd127}: color_data = 12'h333;
			{8'd148, 8'd128}: color_data = 12'h888;
			{8'd148, 8'd129}: color_data = 12'hddd;
			{8'd148, 8'd130}: color_data = 12'heee;
			{8'd148, 8'd131}: color_data = 12'hfff;
			{8'd148, 8'd132}: color_data = 12'hfff;
			{8'd148, 8'd133}: color_data = 12'heee;
			{8'd148, 8'd134}: color_data = 12'hccc;
			{8'd148, 8'd135}: color_data = 12'h777;
			{8'd148, 8'd136}: color_data = 12'h444;
			{8'd149, 8'd102}: color_data = 12'h222;
			{8'd149, 8'd103}: color_data = 12'h222;
			{8'd149, 8'd104}: color_data = 12'h222;
			{8'd149, 8'd105}: color_data = 12'h222;
			{8'd149, 8'd106}: color_data = 12'h222;
			{8'd149, 8'd107}: color_data = 12'h222;
			{8'd149, 8'd108}: color_data = 12'h222;
			{8'd149, 8'd109}: color_data = 12'h222;
			{8'd149, 8'd110}: color_data = 12'h222;
			{8'd149, 8'd111}: color_data = 12'h222;
			{8'd149, 8'd112}: color_data = 12'h222;
			{8'd149, 8'd113}: color_data = 12'h222;
			{8'd149, 8'd114}: color_data = 12'h222;
			{8'd149, 8'd115}: color_data = 12'h222;
			{8'd149, 8'd116}: color_data = 12'h222;
			{8'd149, 8'd117}: color_data = 12'h222;
			{8'd149, 8'd118}: color_data = 12'h111;
			{8'd149, 8'd119}: color_data = 12'h111;
			{8'd149, 8'd120}: color_data = 12'h111;
			{8'd149, 8'd121}: color_data = 12'h111;
			{8'd149, 8'd122}: color_data = 12'h111;
			{8'd149, 8'd123}: color_data = 12'h111;
			{8'd149, 8'd124}: color_data = 12'h111;
			{8'd149, 8'd125}: color_data = 12'h111;
			{8'd149, 8'd126}: color_data = 12'h111;
			{8'd149, 8'd127}: color_data = 12'h111;
			{8'd149, 8'd128}: color_data = 12'h555;
			{8'd149, 8'd129}: color_data = 12'h999;
			{8'd149, 8'd130}: color_data = 12'hccc;
			{8'd149, 8'd131}: color_data = 12'hddd;
			{8'd149, 8'd132}: color_data = 12'hddd;
			{8'd149, 8'd133}: color_data = 12'hccc;
			{8'd149, 8'd134}: color_data = 12'h888;
			{8'd149, 8'd135}: color_data = 12'h444;
			{8'd149, 8'd136}: color_data = 12'h222;
			{8'd150, 8'd107}: color_data = 12'h000;
			{8'd150, 8'd108}: color_data = 12'h222;
			{8'd150, 8'd109}: color_data = 12'h222;
			{8'd150, 8'd110}: color_data = 12'h222;
			{8'd150, 8'd111}: color_data = 12'h222;
			{8'd150, 8'd112}: color_data = 12'h222;
			{8'd150, 8'd113}: color_data = 12'h222;
			{8'd150, 8'd114}: color_data = 12'h222;
			{8'd150, 8'd115}: color_data = 12'h222;
			{8'd150, 8'd116}: color_data = 12'h222;
			{8'd150, 8'd117}: color_data = 12'h111;
			{8'd150, 8'd118}: color_data = 12'h111;
			{8'd150, 8'd119}: color_data = 12'h111;
			{8'd150, 8'd120}: color_data = 12'h111;
			{8'd150, 8'd121}: color_data = 12'h111;
			{8'd150, 8'd122}: color_data = 12'h111;
			{8'd150, 8'd123}: color_data = 12'h111;
			{8'd150, 8'd124}: color_data = 12'h111;
			{8'd150, 8'd125}: color_data = 12'h111;
			{8'd150, 8'd126}: color_data = 12'h111;
			{8'd150, 8'd127}: color_data = 12'h111;
			{8'd150, 8'd128}: color_data = 12'h222;
			{8'd150, 8'd129}: color_data = 12'h555;
			{8'd150, 8'd130}: color_data = 12'h888;
			{8'd150, 8'd131}: color_data = 12'haaa;
			{8'd150, 8'd132}: color_data = 12'haaa;
			{8'd150, 8'd133}: color_data = 12'h888;
			{8'd150, 8'd134}: color_data = 12'h555;
			{8'd150, 8'd135}: color_data = 12'h333;
			{8'd151, 8'd112}: color_data = 12'h000;
			{8'd151, 8'd113}: color_data = 12'h333;
			{8'd151, 8'd114}: color_data = 12'h222;
			{8'd151, 8'd115}: color_data = 12'h111;
			{8'd151, 8'd116}: color_data = 12'h111;
			{8'd151, 8'd117}: color_data = 12'h111;
			{8'd151, 8'd118}: color_data = 12'h111;
			{8'd151, 8'd119}: color_data = 12'h111;
			{8'd151, 8'd120}: color_data = 12'h111;
			{8'd151, 8'd121}: color_data = 12'h111;
			{8'd151, 8'd122}: color_data = 12'h111;
			{8'd151, 8'd123}: color_data = 12'h111;
			{8'd151, 8'd124}: color_data = 12'h111;
			{8'd151, 8'd125}: color_data = 12'h111;
			{8'd151, 8'd126}: color_data = 12'h111;
			{8'd151, 8'd127}: color_data = 12'h111;
			{8'd151, 8'd128}: color_data = 12'h111;
			{8'd151, 8'd129}: color_data = 12'h222;
			{8'd151, 8'd130}: color_data = 12'h444;
			{8'd151, 8'd131}: color_data = 12'h666;
			{8'd151, 8'd132}: color_data = 12'h666;
			{8'd151, 8'd133}: color_data = 12'h555;
			{8'd151, 8'd134}: color_data = 12'h333;
			{8'd152, 8'd34}: color_data = 12'ha11;
			{8'd152, 8'd35}: color_data = 12'ha10;
			{8'd152, 8'd36}: color_data = 12'h700;
			{8'd152, 8'd118}: color_data = 12'h333;
			{8'd152, 8'd119}: color_data = 12'h111;
			{8'd152, 8'd120}: color_data = 12'h111;
			{8'd152, 8'd121}: color_data = 12'h111;
			{8'd152, 8'd122}: color_data = 12'h111;
			{8'd152, 8'd123}: color_data = 12'h111;
			{8'd152, 8'd124}: color_data = 12'h111;
			{8'd152, 8'd125}: color_data = 12'h111;
			{8'd152, 8'd126}: color_data = 12'h111;
			{8'd152, 8'd127}: color_data = 12'h111;
			{8'd152, 8'd128}: color_data = 12'h111;
			{8'd152, 8'd129}: color_data = 12'h222;
			{8'd152, 8'd130}: color_data = 12'h222;
			{8'd152, 8'd131}: color_data = 12'h333;
			{8'd152, 8'd132}: color_data = 12'h333;
			{8'd152, 8'd133}: color_data = 12'h222;
			{8'd153, 8'd33}: color_data = 12'ha01;
			{8'd153, 8'd34}: color_data = 12'hc11;
			{8'd153, 8'd35}: color_data = 12'hc21;
			{8'd153, 8'd36}: color_data = 12'hc21;
			{8'd153, 8'd37}: color_data = 12'hb21;
			{8'd153, 8'd38}: color_data = 12'h920;
			{8'd153, 8'd39}: color_data = 12'h410;
			{8'd153, 8'd40}: color_data = 12'h700;
			{8'd153, 8'd124}: color_data = 12'h111;
			{8'd153, 8'd125}: color_data = 12'h111;
			{8'd153, 8'd126}: color_data = 12'h000;
			{8'd153, 8'd127}: color_data = 12'h000;
			{8'd153, 8'd128}: color_data = 12'h000;
			{8'd153, 8'd129}: color_data = 12'h111;
			{8'd153, 8'd130}: color_data = 12'h222;
			{8'd153, 8'd131}: color_data = 12'h222;
			{8'd153, 8'd132}: color_data = 12'h222;
			{8'd154, 8'd32}: color_data = 12'ha01;
			{8'd154, 8'd33}: color_data = 12'hb11;
			{8'd154, 8'd34}: color_data = 12'hd11;
			{8'd154, 8'd35}: color_data = 12'he21;
			{8'd154, 8'd36}: color_data = 12'hd31;
			{8'd154, 8'd37}: color_data = 12'hc31;
			{8'd154, 8'd38}: color_data = 12'hb31;
			{8'd154, 8'd39}: color_data = 12'ha30;
			{8'd154, 8'd40}: color_data = 12'h820;
			{8'd154, 8'd41}: color_data = 12'h000;
			{8'd154, 8'd129}: color_data = 12'h111;
			{8'd154, 8'd130}: color_data = 12'h222;
			{8'd154, 8'd131}: color_data = 12'h222;
			{8'd154, 8'd132}: color_data = 12'h222;
			{8'd155, 8'd31}: color_data = 12'h000;
			{8'd155, 8'd32}: color_data = 12'ha01;
			{8'd155, 8'd33}: color_data = 12'hd11;
			{8'd155, 8'd34}: color_data = 12'hd11;
			{8'd155, 8'd35}: color_data = 12'hd21;
			{8'd155, 8'd36}: color_data = 12'hd31;
			{8'd155, 8'd37}: color_data = 12'hd31;
			{8'd155, 8'd38}: color_data = 12'he41;
			{8'd155, 8'd39}: color_data = 12'hd41;
			{8'd155, 8'd40}: color_data = 12'hc31;
			{8'd155, 8'd41}: color_data = 12'hc41;
			{8'd155, 8'd42}: color_data = 12'ha40;
			{8'd155, 8'd43}: color_data = 12'h930;
			{8'd155, 8'd44}: color_data = 12'h550;
			{8'd156, 8'd30}: color_data = 12'h700;
			{8'd156, 8'd31}: color_data = 12'ha01;
			{8'd156, 8'd32}: color_data = 12'hc01;
			{8'd156, 8'd33}: color_data = 12'hd11;
			{8'd156, 8'd34}: color_data = 12'hd11;
			{8'd156, 8'd35}: color_data = 12'hd21;
			{8'd156, 8'd36}: color_data = 12'hd31;
			{8'd156, 8'd37}: color_data = 12'hd31;
			{8'd156, 8'd38}: color_data = 12'hd31;
			{8'd156, 8'd39}: color_data = 12'he41;
			{8'd156, 8'd40}: color_data = 12'he41;
			{8'd156, 8'd41}: color_data = 12'he51;
			{8'd156, 8'd42}: color_data = 12'hd51;
			{8'd156, 8'd43}: color_data = 12'hc51;
			{8'd156, 8'd44}: color_data = 12'hb50;
			{8'd156, 8'd45}: color_data = 12'ha50;
			{8'd156, 8'd46}: color_data = 12'h841;
			{8'd156, 8'd47}: color_data = 12'h940;
			{8'd157, 8'd30}: color_data = 12'h901;
			{8'd157, 8'd31}: color_data = 12'hb01;
			{8'd157, 8'd32}: color_data = 12'hd01;
			{8'd157, 8'd33}: color_data = 12'hd11;
			{8'd157, 8'd34}: color_data = 12'hd11;
			{8'd157, 8'd35}: color_data = 12'hd21;
			{8'd157, 8'd36}: color_data = 12'hd31;
			{8'd157, 8'd37}: color_data = 12'hd31;
			{8'd157, 8'd38}: color_data = 12'hd31;
			{8'd157, 8'd39}: color_data = 12'he41;
			{8'd157, 8'd40}: color_data = 12'he41;
			{8'd157, 8'd41}: color_data = 12'he51;
			{8'd157, 8'd42}: color_data = 12'he51;
			{8'd157, 8'd43}: color_data = 12'he61;
			{8'd157, 8'd44}: color_data = 12'hd61;
			{8'd157, 8'd45}: color_data = 12'hd61;
			{8'd157, 8'd46}: color_data = 12'hb51;
			{8'd157, 8'd47}: color_data = 12'ha51;
			{8'd157, 8'd48}: color_data = 12'ha60;
			{8'd157, 8'd49}: color_data = 12'ha51;
			{8'd158, 8'd30}: color_data = 12'ha01;
			{8'd158, 8'd31}: color_data = 12'hc01;
			{8'd158, 8'd32}: color_data = 12'hd01;
			{8'd158, 8'd33}: color_data = 12'hd11;
			{8'd158, 8'd34}: color_data = 12'hd11;
			{8'd158, 8'd35}: color_data = 12'hd21;
			{8'd158, 8'd36}: color_data = 12'hd31;
			{8'd158, 8'd37}: color_data = 12'hd31;
			{8'd158, 8'd38}: color_data = 12'hd31;
			{8'd158, 8'd39}: color_data = 12'he41;
			{8'd158, 8'd40}: color_data = 12'he41;
			{8'd158, 8'd41}: color_data = 12'he51;
			{8'd158, 8'd42}: color_data = 12'he51;
			{8'd158, 8'd43}: color_data = 12'he51;
			{8'd158, 8'd44}: color_data = 12'he61;
			{8'd158, 8'd45}: color_data = 12'he71;
			{8'd158, 8'd46}: color_data = 12'he71;
			{8'd158, 8'd47}: color_data = 12'hd71;
			{8'd158, 8'd48}: color_data = 12'hc61;
			{8'd158, 8'd49}: color_data = 12'hb60;
			{8'd158, 8'd50}: color_data = 12'hb60;
			{8'd158, 8'd51}: color_data = 12'ha50;
			{8'd158, 8'd52}: color_data = 12'h000;
			{8'd159, 8'd30}: color_data = 12'hb01;
			{8'd159, 8'd31}: color_data = 12'hc01;
			{8'd159, 8'd32}: color_data = 12'he01;
			{8'd159, 8'd33}: color_data = 12'hd11;
			{8'd159, 8'd34}: color_data = 12'he21;
			{8'd159, 8'd35}: color_data = 12'he21;
			{8'd159, 8'd36}: color_data = 12'he31;
			{8'd159, 8'd37}: color_data = 12'he31;
			{8'd159, 8'd38}: color_data = 12'he41;
			{8'd159, 8'd39}: color_data = 12'he41;
			{8'd159, 8'd40}: color_data = 12'he41;
			{8'd159, 8'd41}: color_data = 12'he51;
			{8'd159, 8'd42}: color_data = 12'he51;
			{8'd159, 8'd43}: color_data = 12'he61;
			{8'd159, 8'd44}: color_data = 12'he61;
			{8'd159, 8'd45}: color_data = 12'he61;
			{8'd159, 8'd46}: color_data = 12'he71;
			{8'd159, 8'd47}: color_data = 12'he71;
			{8'd159, 8'd48}: color_data = 12'he71;
			{8'd159, 8'd49}: color_data = 12'hd70;
			{8'd159, 8'd50}: color_data = 12'hd70;
			{8'd159, 8'd51}: color_data = 12'hc70;
			{8'd159, 8'd52}: color_data = 12'hb70;
			{8'd159, 8'd53}: color_data = 12'h960;
			{8'd159, 8'd54}: color_data = 12'h850;
			{8'd160, 8'd30}: color_data = 12'hb01;
			{8'd160, 8'd31}: color_data = 12'hc01;
			{8'd160, 8'd32}: color_data = 12'hc01;
			{8'd160, 8'd33}: color_data = 12'hd01;
			{8'd160, 8'd34}: color_data = 12'hd11;
			{8'd160, 8'd35}: color_data = 12'hd21;
			{8'd160, 8'd36}: color_data = 12'hd31;
			{8'd160, 8'd37}: color_data = 12'hd31;
			{8'd160, 8'd38}: color_data = 12'hd31;
			{8'd160, 8'd39}: color_data = 12'he41;
			{8'd160, 8'd40}: color_data = 12'he41;
			{8'd160, 8'd41}: color_data = 12'he51;
			{8'd160, 8'd42}: color_data = 12'he51;
			{8'd160, 8'd43}: color_data = 12'he51;
			{8'd160, 8'd44}: color_data = 12'hd61;
			{8'd160, 8'd45}: color_data = 12'hc61;
			{8'd160, 8'd46}: color_data = 12'he71;
			{8'd160, 8'd47}: color_data = 12'he71;
			{8'd160, 8'd48}: color_data = 12'he71;
			{8'd160, 8'd49}: color_data = 12'he80;
			{8'd160, 8'd50}: color_data = 12'he80;
			{8'd160, 8'd51}: color_data = 12'he80;
			{8'd160, 8'd52}: color_data = 12'he80;
			{8'd160, 8'd53}: color_data = 12'hc80;
			{8'd160, 8'd54}: color_data = 12'hb70;
			{8'd160, 8'd55}: color_data = 12'hb70;
			{8'd161, 8'd45}: color_data = 12'hb51;
			{8'd161, 8'd46}: color_data = 12'hd61;
			{8'd161, 8'd47}: color_data = 12'he71;
			{8'd161, 8'd48}: color_data = 12'he71;
			{8'd161, 8'd49}: color_data = 12'he80;
			{8'd161, 8'd50}: color_data = 12'he80;
			{8'd161, 8'd51}: color_data = 12'he80;
			{8'd161, 8'd52}: color_data = 12'he80;
			{8'd161, 8'd53}: color_data = 12'he90;
			{8'd161, 8'd54}: color_data = 12'he90;
			{8'd161, 8'd55}: color_data = 12'hc80;
			{8'd161, 8'd56}: color_data = 12'h770;
			{8'd162, 8'd45}: color_data = 12'hd61;
			{8'd162, 8'd46}: color_data = 12'hd61;
			{8'd162, 8'd47}: color_data = 12'he71;
			{8'd162, 8'd48}: color_data = 12'he71;
			{8'd162, 8'd49}: color_data = 12'he80;
			{8'd162, 8'd50}: color_data = 12'he80;
			{8'd162, 8'd51}: color_data = 12'he80;
			{8'd162, 8'd52}: color_data = 12'he80;
			{8'd162, 8'd53}: color_data = 12'he90;
			{8'd162, 8'd54}: color_data = 12'hd90;
			{8'd162, 8'd55}: color_data = 12'hb80;
			{8'd162, 8'd56}: color_data = 12'hb70;
			{8'd163, 8'd45}: color_data = 12'he61;
			{8'd163, 8'd46}: color_data = 12'he61;
			{8'd163, 8'd47}: color_data = 12'he71;
			{8'd163, 8'd48}: color_data = 12'he71;
			{8'd163, 8'd49}: color_data = 12'he80;
			{8'd163, 8'd50}: color_data = 12'he80;
			{8'd163, 8'd51}: color_data = 12'he80;
			{8'd163, 8'd52}: color_data = 12'he80;
			{8'd163, 8'd53}: color_data = 12'he90;
			{8'd163, 8'd54}: color_data = 12'hd90;
			{8'd163, 8'd55}: color_data = 12'hb80;
			{8'd163, 8'd56}: color_data = 12'hf00;
			{8'd164, 8'd45}: color_data = 12'hc61;
			{8'd164, 8'd46}: color_data = 12'hd61;
			{8'd164, 8'd47}: color_data = 12'he71;
			{8'd164, 8'd48}: color_data = 12'he71;
			{8'd164, 8'd49}: color_data = 12'he80;
			{8'd164, 8'd50}: color_data = 12'he80;
			{8'd164, 8'd51}: color_data = 12'he80;
			{8'd164, 8'd52}: color_data = 12'hd80;
			{8'd164, 8'd53}: color_data = 12'hd80;
			{8'd164, 8'd54}: color_data = 12'hc80;
			{8'd164, 8'd55}: color_data = 12'hb70;
			{8'd165, 8'd33}: color_data = 12'h000;
			{8'd165, 8'd34}: color_data = 12'h000;
			{8'd165, 8'd35}: color_data = 12'h710;
			{8'd165, 8'd36}: color_data = 12'h810;
			{8'd165, 8'd37}: color_data = 12'h710;
			{8'd165, 8'd38}: color_data = 12'h710;
			{8'd165, 8'd39}: color_data = 12'h820;
			{8'd165, 8'd40}: color_data = 12'h820;
			{8'd165, 8'd41}: color_data = 12'h820;
			{8'd165, 8'd42}: color_data = 12'h830;
			{8'd165, 8'd43}: color_data = 12'h830;
			{8'd165, 8'd44}: color_data = 12'h830;
			{8'd165, 8'd45}: color_data = 12'h940;
			{8'd165, 8'd46}: color_data = 12'hd61;
			{8'd165, 8'd47}: color_data = 12'he71;
			{8'd165, 8'd48}: color_data = 12'he71;
			{8'd165, 8'd49}: color_data = 12'he80;
			{8'd165, 8'd50}: color_data = 12'hd80;
			{8'd165, 8'd51}: color_data = 12'hc70;
			{8'd165, 8'd52}: color_data = 12'hc70;
			{8'd165, 8'd53}: color_data = 12'hb70;
			{8'd166, 8'd32}: color_data = 12'hb10;
			{8'd166, 8'd33}: color_data = 12'ha11;
			{8'd166, 8'd34}: color_data = 12'ha11;
			{8'd166, 8'd35}: color_data = 12'h911;
			{8'd166, 8'd36}: color_data = 12'h920;
			{8'd166, 8'd37}: color_data = 12'h920;
			{8'd166, 8'd38}: color_data = 12'h920;
			{8'd166, 8'd39}: color_data = 12'h930;
			{8'd166, 8'd40}: color_data = 12'ha30;
			{8'd166, 8'd41}: color_data = 12'ha30;
			{8'd166, 8'd42}: color_data = 12'ha40;
			{8'd166, 8'd43}: color_data = 12'ha40;
			{8'd166, 8'd44}: color_data = 12'ha41;
			{8'd166, 8'd45}: color_data = 12'hc51;
			{8'd166, 8'd46}: color_data = 12'he71;
			{8'd166, 8'd47}: color_data = 12'he71;
			{8'd166, 8'd48}: color_data = 12'hd71;
			{8'd166, 8'd49}: color_data = 12'hc60;
			{8'd166, 8'd50}: color_data = 12'hb60;
			{8'd166, 8'd51}: color_data = 12'h950;
			{8'd166, 8'd52}: color_data = 12'h730;
			{8'd167, 8'd32}: color_data = 12'ha11;
			{8'd167, 8'd33}: color_data = 12'hc11;
			{8'd167, 8'd34}: color_data = 12'hd11;
			{8'd167, 8'd35}: color_data = 12'hd21;
			{8'd167, 8'd36}: color_data = 12'hd31;
			{8'd167, 8'd37}: color_data = 12'hd31;
			{8'd167, 8'd38}: color_data = 12'hd31;
			{8'd167, 8'd39}: color_data = 12'hd41;
			{8'd167, 8'd40}: color_data = 12'hd41;
			{8'd167, 8'd41}: color_data = 12'hd51;
			{8'd167, 8'd42}: color_data = 12'he51;
			{8'd167, 8'd43}: color_data = 12'he51;
			{8'd167, 8'd44}: color_data = 12'he61;
			{8'd167, 8'd45}: color_data = 12'he61;
			{8'd167, 8'd46}: color_data = 12'hd61;
			{8'd167, 8'd47}: color_data = 12'hb60;
			{8'd167, 8'd48}: color_data = 12'ha50;
			{8'd167, 8'd49}: color_data = 12'h840;
			{8'd168, 8'd32}: color_data = 12'h900;
			{8'd168, 8'd33}: color_data = 12'hb11;
			{8'd168, 8'd34}: color_data = 12'hd11;
			{8'd168, 8'd35}: color_data = 12'hd21;
			{8'd168, 8'd36}: color_data = 12'hd31;
			{8'd168, 8'd37}: color_data = 12'hd31;
			{8'd168, 8'd38}: color_data = 12'hd41;
			{8'd168, 8'd39}: color_data = 12'he41;
			{8'd168, 8'd40}: color_data = 12'he41;
			{8'd168, 8'd41}: color_data = 12'he51;
			{8'd168, 8'd42}: color_data = 12'he51;
			{8'd168, 8'd43}: color_data = 12'he61;
			{8'd168, 8'd44}: color_data = 12'hc51;
			{8'd168, 8'd45}: color_data = 12'hc50;
			{8'd168, 8'd46}: color_data = 12'ha50;
			{8'd168, 8'd47}: color_data = 12'h840;
			{8'd168, 8'd48}: color_data = 12'h741;
			{8'd169, 8'd33}: color_data = 12'ha10;
			{8'd169, 8'd34}: color_data = 12'hb11;
			{8'd169, 8'd35}: color_data = 12'hd21;
			{8'd169, 8'd36}: color_data = 12'hd31;
			{8'd169, 8'd37}: color_data = 12'hd31;
			{8'd169, 8'd38}: color_data = 12'hd31;
			{8'd169, 8'd39}: color_data = 12'he41;
			{8'd169, 8'd40}: color_data = 12'he41;
			{8'd169, 8'd41}: color_data = 12'hd51;
			{8'd169, 8'd42}: color_data = 12'hc41;
			{8'd169, 8'd43}: color_data = 12'hb41;
			{8'd169, 8'd44}: color_data = 12'ha40;
			{8'd169, 8'd45}: color_data = 12'ha31;
			{8'd170, 8'd34}: color_data = 12'ha11;
			{8'd170, 8'd35}: color_data = 12'hc21;
			{8'd170, 8'd36}: color_data = 12'he31;
			{8'd170, 8'd37}: color_data = 12'hd31;
			{8'd170, 8'd38}: color_data = 12'hd31;
			{8'd170, 8'd39}: color_data = 12'hd41;
			{8'd170, 8'd40}: color_data = 12'hb30;
			{8'd170, 8'd41}: color_data = 12'hb30;
			{8'd170, 8'd42}: color_data = 12'ha41;
			{8'd170, 8'd43}: color_data = 12'ha50;
			{8'd171, 8'd35}: color_data = 12'ha21;
			{8'd171, 8'd36}: color_data = 12'hc21;
			{8'd171, 8'd37}: color_data = 12'hd31;
			{8'd171, 8'd38}: color_data = 12'hc31;
			{8'd171, 8'd39}: color_data = 12'ha30;
			{8'd171, 8'd40}: color_data = 12'h920;
			{8'd171, 8'd41}: color_data = 12'h610;
			{8'd172, 8'd35}: color_data = 12'h910;
			{8'd172, 8'd36}: color_data = 12'ha21;
			{8'd172, 8'd37}: color_data = 12'hb31;
			{8'd172, 8'd38}: color_data = 12'hc31;
			{8'd176, 8'd34}: color_data = 12'h720;
			{8'd176, 8'd35}: color_data = 12'h820;
			{8'd176, 8'd36}: color_data = 12'h720;
			{8'd176, 8'd37}: color_data = 12'h000;
			{8'd177, 8'd33}: color_data = 12'h921;
			{8'd177, 8'd34}: color_data = 12'ha21;
			{8'd177, 8'd35}: color_data = 12'ha20;
			{8'd177, 8'd36}: color_data = 12'ha20;
			{8'd177, 8'd37}: color_data = 12'ha30;
			{8'd177, 8'd38}: color_data = 12'h930;
			{8'd178, 8'd33}: color_data = 12'ha21;
			{8'd178, 8'd34}: color_data = 12'hc31;
			{8'd178, 8'd35}: color_data = 12'hd31;
			{8'd178, 8'd36}: color_data = 12'hd41;
			{8'd178, 8'd37}: color_data = 12'hd41;
			{8'd178, 8'd38}: color_data = 12'hb41;
			{8'd178, 8'd39}: color_data = 12'ha30;
			{8'd178, 8'd40}: color_data = 12'ha40;
			{8'd178, 8'd41}: color_data = 12'ha40;
			{8'd178, 8'd42}: color_data = 12'ha50;
			{8'd178, 8'd43}: color_data = 12'ha50;
			{8'd178, 8'd44}: color_data = 12'hb50;
			{8'd178, 8'd45}: color_data = 12'hb50;
			{8'd178, 8'd46}: color_data = 12'hb60;
			{8'd178, 8'd47}: color_data = 12'hb60;
			{8'd178, 8'd48}: color_data = 12'hb60;
			{8'd178, 8'd49}: color_data = 12'hb70;
			{8'd178, 8'd50}: color_data = 12'hb70;
			{8'd178, 8'd51}: color_data = 12'hb70;
			{8'd178, 8'd52}: color_data = 12'hb80;
			{8'd178, 8'd53}: color_data = 12'hb71;
			{8'd179, 8'd33}: color_data = 12'hc31;
			{8'd179, 8'd34}: color_data = 12'hd31;
			{8'd179, 8'd35}: color_data = 12'he31;
			{8'd179, 8'd36}: color_data = 12'he41;
			{8'd179, 8'd37}: color_data = 12'he41;
			{8'd179, 8'd38}: color_data = 12'hd51;
			{8'd179, 8'd39}: color_data = 12'hc41;
			{8'd179, 8'd40}: color_data = 12'hc51;
			{8'd179, 8'd41}: color_data = 12'hc51;
			{8'd179, 8'd42}: color_data = 12'hc61;
			{8'd179, 8'd43}: color_data = 12'hc61;
			{8'd179, 8'd44}: color_data = 12'hc61;
			{8'd179, 8'd45}: color_data = 12'hc70;
			{8'd179, 8'd46}: color_data = 12'hc70;
			{8'd179, 8'd47}: color_data = 12'hd70;
			{8'd179, 8'd48}: color_data = 12'hd80;
			{8'd179, 8'd49}: color_data = 12'hd80;
			{8'd179, 8'd50}: color_data = 12'hd80;
			{8'd179, 8'd51}: color_data = 12'hd90;
			{8'd179, 8'd52}: color_data = 12'hd90;
			{8'd179, 8'd53}: color_data = 12'hc80;
			{8'd180, 8'd33}: color_data = 12'hd31;
			{8'd180, 8'd34}: color_data = 12'hd31;
			{8'd180, 8'd35}: color_data = 12'he31;
			{8'd180, 8'd36}: color_data = 12'he41;
			{8'd180, 8'd37}: color_data = 12'he41;
			{8'd180, 8'd38}: color_data = 12'he51;
			{8'd180, 8'd39}: color_data = 12'he51;
			{8'd180, 8'd40}: color_data = 12'he61;
			{8'd180, 8'd41}: color_data = 12'he61;
			{8'd180, 8'd42}: color_data = 12'he61;
			{8'd180, 8'd43}: color_data = 12'he71;
			{8'd180, 8'd44}: color_data = 12'he71;
			{8'd180, 8'd45}: color_data = 12'he81;
			{8'd180, 8'd46}: color_data = 12'he80;
			{8'd180, 8'd47}: color_data = 12'he80;
			{8'd180, 8'd48}: color_data = 12'he80;
			{8'd180, 8'd49}: color_data = 12'he90;
			{8'd180, 8'd50}: color_data = 12'he90;
			{8'd180, 8'd51}: color_data = 12'he90;
			{8'd180, 8'd52}: color_data = 12'hea0;
			{8'd180, 8'd53}: color_data = 12'hd90;
			{8'd181, 8'd33}: color_data = 12'hd31;
			{8'd181, 8'd34}: color_data = 12'hd31;
			{8'd181, 8'd35}: color_data = 12'he31;
			{8'd181, 8'd36}: color_data = 12'he41;
			{8'd181, 8'd37}: color_data = 12'he41;
			{8'd181, 8'd38}: color_data = 12'he51;
			{8'd181, 8'd39}: color_data = 12'he51;
			{8'd181, 8'd40}: color_data = 12'he61;
			{8'd181, 8'd41}: color_data = 12'he61;
			{8'd181, 8'd42}: color_data = 12'he61;
			{8'd181, 8'd43}: color_data = 12'he71;
			{8'd181, 8'd44}: color_data = 12'he71;
			{8'd181, 8'd45}: color_data = 12'he71;
			{8'd181, 8'd46}: color_data = 12'he80;
			{8'd181, 8'd47}: color_data = 12'he80;
			{8'd181, 8'd48}: color_data = 12'he80;
			{8'd181, 8'd49}: color_data = 12'he90;
			{8'd181, 8'd50}: color_data = 12'he90;
			{8'd181, 8'd51}: color_data = 12'he90;
			{8'd181, 8'd52}: color_data = 12'hea0;
			{8'd181, 8'd53}: color_data = 12'hd90;
			{8'd182, 8'd33}: color_data = 12'hc31;
			{8'd182, 8'd34}: color_data = 12'hd31;
			{8'd182, 8'd35}: color_data = 12'he31;
			{8'd182, 8'd36}: color_data = 12'he41;
			{8'd182, 8'd37}: color_data = 12'he41;
			{8'd182, 8'd38}: color_data = 12'he51;
			{8'd182, 8'd39}: color_data = 12'he51;
			{8'd182, 8'd40}: color_data = 12'he61;
			{8'd182, 8'd41}: color_data = 12'he61;
			{8'd182, 8'd42}: color_data = 12'he61;
			{8'd182, 8'd43}: color_data = 12'he71;
			{8'd182, 8'd44}: color_data = 12'he71;
			{8'd182, 8'd45}: color_data = 12'he71;
			{8'd182, 8'd46}: color_data = 12'he80;
			{8'd182, 8'd47}: color_data = 12'he80;
			{8'd182, 8'd48}: color_data = 12'he80;
			{8'd182, 8'd49}: color_data = 12'he90;
			{8'd182, 8'd50}: color_data = 12'he90;
			{8'd182, 8'd51}: color_data = 12'he90;
			{8'd182, 8'd52}: color_data = 12'hea0;
			{8'd182, 8'd53}: color_data = 12'hd90;
			{8'd183, 8'd33}: color_data = 12'hc21;
			{8'd183, 8'd34}: color_data = 12'hd31;
			{8'd183, 8'd35}: color_data = 12'he31;
			{8'd183, 8'd36}: color_data = 12'he41;
			{8'd183, 8'd37}: color_data = 12'he41;
			{8'd183, 8'd38}: color_data = 12'he51;
			{8'd183, 8'd39}: color_data = 12'he51;
			{8'd183, 8'd40}: color_data = 12'he61;
			{8'd183, 8'd41}: color_data = 12'he61;
			{8'd183, 8'd42}: color_data = 12'he61;
			{8'd183, 8'd43}: color_data = 12'he71;
			{8'd183, 8'd44}: color_data = 12'he71;
			{8'd183, 8'd45}: color_data = 12'he71;
			{8'd183, 8'd46}: color_data = 12'he80;
			{8'd183, 8'd47}: color_data = 12'he80;
			{8'd183, 8'd48}: color_data = 12'he80;
			{8'd183, 8'd49}: color_data = 12'he90;
			{8'd183, 8'd50}: color_data = 12'he90;
			{8'd183, 8'd51}: color_data = 12'he90;
			{8'd183, 8'd52}: color_data = 12'hea0;
			{8'd183, 8'd53}: color_data = 12'hd90;
			{8'd184, 8'd33}: color_data = 12'hc21;
			{8'd184, 8'd34}: color_data = 12'hd31;
			{8'd184, 8'd35}: color_data = 12'he31;
			{8'd184, 8'd36}: color_data = 12'he41;
			{8'd184, 8'd37}: color_data = 12'he41;
			{8'd184, 8'd38}: color_data = 12'he51;
			{8'd184, 8'd39}: color_data = 12'he51;
			{8'd184, 8'd40}: color_data = 12'he61;
			{8'd184, 8'd41}: color_data = 12'he61;
			{8'd184, 8'd42}: color_data = 12'he61;
			{8'd184, 8'd43}: color_data = 12'he71;
			{8'd184, 8'd44}: color_data = 12'he71;
			{8'd184, 8'd45}: color_data = 12'hd71;
			{8'd184, 8'd46}: color_data = 12'hc70;
			{8'd184, 8'd47}: color_data = 12'hd80;
			{8'd184, 8'd48}: color_data = 12'he80;
			{8'd184, 8'd49}: color_data = 12'he90;
			{8'd184, 8'd50}: color_data = 12'he90;
			{8'd184, 8'd51}: color_data = 12'he90;
			{8'd184, 8'd52}: color_data = 12'hea0;
			{8'd184, 8'd53}: color_data = 12'hd90;
			{8'd185, 8'd33}: color_data = 12'hc21;
			{8'd185, 8'd34}: color_data = 12'hd31;
			{8'd185, 8'd35}: color_data = 12'hd31;
			{8'd185, 8'd36}: color_data = 12'hd41;
			{8'd185, 8'd37}: color_data = 12'he41;
			{8'd185, 8'd38}: color_data = 12'hd51;
			{8'd185, 8'd39}: color_data = 12'hc41;
			{8'd185, 8'd40}: color_data = 12'hd51;
			{8'd185, 8'd41}: color_data = 12'he61;
			{8'd185, 8'd42}: color_data = 12'he61;
			{8'd185, 8'd43}: color_data = 12'he71;
			{8'd185, 8'd44}: color_data = 12'he71;
			{8'd185, 8'd45}: color_data = 12'hb60;
			{8'd185, 8'd46}: color_data = 12'h840;
			{8'd185, 8'd47}: color_data = 12'hb60;
			{8'd185, 8'd48}: color_data = 12'he80;
			{8'd185, 8'd49}: color_data = 12'he90;
			{8'd185, 8'd50}: color_data = 12'he90;
			{8'd185, 8'd51}: color_data = 12'he90;
			{8'd185, 8'd52}: color_data = 12'hea0;
			{8'd185, 8'd53}: color_data = 12'hd90;
			{8'd186, 8'd33}: color_data = 12'hb21;
			{8'd186, 8'd34}: color_data = 12'hd31;
			{8'd186, 8'd35}: color_data = 12'hd31;
			{8'd186, 8'd36}: color_data = 12'hd41;
			{8'd186, 8'd37}: color_data = 12'he41;
			{8'd186, 8'd38}: color_data = 12'hb40;
			{8'd186, 8'd39}: color_data = 12'h720;
			{8'd186, 8'd40}: color_data = 12'hc51;
			{8'd186, 8'd41}: color_data = 12'he61;
			{8'd186, 8'd42}: color_data = 12'he61;
			{8'd186, 8'd43}: color_data = 12'he71;
			{8'd186, 8'd44}: color_data = 12'he71;
			{8'd186, 8'd45}: color_data = 12'hc60;
			{8'd186, 8'd46}: color_data = 12'h730;
			{8'd186, 8'd47}: color_data = 12'hc70;
			{8'd186, 8'd48}: color_data = 12'he80;
			{8'd186, 8'd49}: color_data = 12'he90;
			{8'd186, 8'd50}: color_data = 12'he90;
			{8'd186, 8'd51}: color_data = 12'he90;
			{8'd186, 8'd52}: color_data = 12'he90;
			{8'd186, 8'd53}: color_data = 12'hd90;
			{8'd187, 8'd32}: color_data = 12'hc11;
			{8'd187, 8'd33}: color_data = 12'hc21;
			{8'd187, 8'd34}: color_data = 12'hd31;
			{8'd187, 8'd35}: color_data = 12'hd31;
			{8'd187, 8'd36}: color_data = 12'hd41;
			{8'd187, 8'd37}: color_data = 12'he41;
			{8'd187, 8'd38}: color_data = 12'hb40;
			{8'd187, 8'd39}: color_data = 12'h310;
			{8'd187, 8'd40}: color_data = 12'hd51;
			{8'd187, 8'd41}: color_data = 12'he61;
			{8'd187, 8'd42}: color_data = 12'he61;
			{8'd187, 8'd43}: color_data = 12'he71;
			{8'd187, 8'd44}: color_data = 12'he71;
			{8'd187, 8'd45}: color_data = 12'hd71;
			{8'd187, 8'd46}: color_data = 12'hb60;
			{8'd187, 8'd47}: color_data = 12'hc70;
			{8'd187, 8'd48}: color_data = 12'he80;
			{8'd187, 8'd49}: color_data = 12'he90;
			{8'd187, 8'd50}: color_data = 12'he90;
			{8'd187, 8'd51}: color_data = 12'he90;
			{8'd187, 8'd52}: color_data = 12'hd90;
			{8'd187, 8'd53}: color_data = 12'hd80;
			{8'd188, 8'd32}: color_data = 12'hb21;
			{8'd188, 8'd33}: color_data = 12'hc21;
			{8'd188, 8'd34}: color_data = 12'he31;
			{8'd188, 8'd35}: color_data = 12'hd31;
			{8'd188, 8'd36}: color_data = 12'hd41;
			{8'd188, 8'd37}: color_data = 12'he41;
			{8'd188, 8'd38}: color_data = 12'hb40;
			{8'd188, 8'd40}: color_data = 12'he61;
			{8'd188, 8'd41}: color_data = 12'he61;
			{8'd188, 8'd42}: color_data = 12'he61;
			{8'd188, 8'd43}: color_data = 12'he71;
			{8'd188, 8'd44}: color_data = 12'he71;
			{8'd188, 8'd45}: color_data = 12'hd70;
			{8'd188, 8'd46}: color_data = 12'hb70;
			{8'd188, 8'd47}: color_data = 12'hc70;
			{8'd188, 8'd48}: color_data = 12'he80;
			{8'd188, 8'd49}: color_data = 12'he90;
			{8'd188, 8'd50}: color_data = 12'he90;
			{8'd188, 8'd51}: color_data = 12'he90;
			{8'd188, 8'd52}: color_data = 12'hd90;
			{8'd188, 8'd53}: color_data = 12'hc80;
			{8'd189, 8'd32}: color_data = 12'hc21;
			{8'd189, 8'd33}: color_data = 12'hd21;
			{8'd189, 8'd34}: color_data = 12'hd31;
			{8'd189, 8'd35}: color_data = 12'hd31;
			{8'd189, 8'd36}: color_data = 12'hd41;
			{8'd189, 8'd37}: color_data = 12'he41;
			{8'd189, 8'd38}: color_data = 12'hb30;
			{8'd189, 8'd39}: color_data = 12'h310;
			{8'd189, 8'd40}: color_data = 12'hd51;
			{8'd189, 8'd41}: color_data = 12'he61;
			{8'd189, 8'd42}: color_data = 12'he61;
			{8'd189, 8'd43}: color_data = 12'he71;
			{8'd189, 8'd44}: color_data = 12'he71;
			{8'd189, 8'd45}: color_data = 12'hd71;
			{8'd189, 8'd46}: color_data = 12'ha70;
			{8'd189, 8'd47}: color_data = 12'hc70;
			{8'd189, 8'd48}: color_data = 12'he80;
			{8'd189, 8'd49}: color_data = 12'he90;
			{8'd189, 8'd50}: color_data = 12'he90;
			{8'd189, 8'd51}: color_data = 12'he90;
			{8'd189, 8'd52}: color_data = 12'hd90;
			{8'd189, 8'd53}: color_data = 12'hc80;
			{8'd190, 8'd32}: color_data = 12'hc21;
			{8'd190, 8'd33}: color_data = 12'hd21;
			{8'd190, 8'd34}: color_data = 12'hd31;
			{8'd190, 8'd35}: color_data = 12'hd31;
			{8'd190, 8'd36}: color_data = 12'hd41;
			{8'd190, 8'd37}: color_data = 12'he41;
			{8'd190, 8'd38}: color_data = 12'hc40;
			{8'd190, 8'd39}: color_data = 12'h510;
			{8'd190, 8'd40}: color_data = 12'hd51;
			{8'd190, 8'd41}: color_data = 12'he61;
			{8'd190, 8'd42}: color_data = 12'he61;
			{8'd190, 8'd43}: color_data = 12'he71;
			{8'd190, 8'd44}: color_data = 12'he71;
			{8'd190, 8'd45}: color_data = 12'hc60;
			{8'd190, 8'd47}: color_data = 12'hd80;
			{8'd190, 8'd48}: color_data = 12'he80;
			{8'd190, 8'd49}: color_data = 12'he90;
			{8'd190, 8'd50}: color_data = 12'he90;
			{8'd190, 8'd51}: color_data = 12'he90;
			{8'd190, 8'd52}: color_data = 12'hd90;
			{8'd190, 8'd53}: color_data = 12'hc80;
			{8'd191, 8'd32}: color_data = 12'hc21;
			{8'd191, 8'd33}: color_data = 12'hd21;
			{8'd191, 8'd34}: color_data = 12'hd31;
			{8'd191, 8'd35}: color_data = 12'hd31;
			{8'd191, 8'd36}: color_data = 12'hd41;
			{8'd191, 8'd37}: color_data = 12'he41;
			{8'd191, 8'd38}: color_data = 12'hd41;
			{8'd191, 8'd39}: color_data = 12'hc41;
			{8'd191, 8'd40}: color_data = 12'hc51;
			{8'd191, 8'd41}: color_data = 12'hd61;
			{8'd191, 8'd42}: color_data = 12'hd61;
			{8'd191, 8'd43}: color_data = 12'hc60;
			{8'd191, 8'd44}: color_data = 12'hb60;
			{8'd191, 8'd45}: color_data = 12'hb50;
			{8'd191, 8'd47}: color_data = 12'he80;
			{8'd191, 8'd48}: color_data = 12'he80;
			{8'd191, 8'd49}: color_data = 12'he90;
			{8'd191, 8'd50}: color_data = 12'he90;
			{8'd191, 8'd51}: color_data = 12'he90;
			{8'd191, 8'd52}: color_data = 12'hd90;
			{8'd191, 8'd53}: color_data = 12'hc80;
			{8'd192, 8'd32}: color_data = 12'hc21;
			{8'd192, 8'd33}: color_data = 12'hd21;
			{8'd192, 8'd34}: color_data = 12'hd31;
			{8'd192, 8'd35}: color_data = 12'hd31;
			{8'd192, 8'd36}: color_data = 12'hd41;
			{8'd192, 8'd37}: color_data = 12'he41;
			{8'd192, 8'd38}: color_data = 12'hd41;
			{8'd192, 8'd39}: color_data = 12'hd40;
			{8'd192, 8'd41}: color_data = 12'hc61;
			{8'd192, 8'd42}: color_data = 12'hd61;
			{8'd192, 8'd43}: color_data = 12'hc51;
			{8'd192, 8'd44}: color_data = 12'h950;
			{8'd192, 8'd45}: color_data = 12'hf00;
			{8'd192, 8'd47}: color_data = 12'hd80;
			{8'd192, 8'd48}: color_data = 12'he80;
			{8'd192, 8'd49}: color_data = 12'he90;
			{8'd192, 8'd50}: color_data = 12'he90;
			{8'd192, 8'd51}: color_data = 12'he90;
			{8'd192, 8'd52}: color_data = 12'hd90;
			{8'd192, 8'd53}: color_data = 12'hc80;
			{8'd193, 8'd31}: color_data = 12'hc21;
			{8'd193, 8'd32}: color_data = 12'hc21;
			{8'd193, 8'd33}: color_data = 12'hd21;
			{8'd193, 8'd34}: color_data = 12'hd31;
			{8'd193, 8'd35}: color_data = 12'hd31;
			{8'd193, 8'd36}: color_data = 12'hd41;
			{8'd193, 8'd37}: color_data = 12'he41;
			{8'd193, 8'd38}: color_data = 12'hd41;
			{8'd193, 8'd39}: color_data = 12'he40;
			{8'd193, 8'd47}: color_data = 12'hc70;
			{8'd193, 8'd48}: color_data = 12'he80;
			{8'd193, 8'd49}: color_data = 12'he90;
			{8'd193, 8'd50}: color_data = 12'he90;
			{8'd193, 8'd51}: color_data = 12'he90;
			{8'd193, 8'd52}: color_data = 12'hd90;
			{8'd193, 8'd53}: color_data = 12'ha70;
			{8'd194, 8'd31}: color_data = 12'hc21;
			{8'd194, 8'd32}: color_data = 12'hc21;
			{8'd194, 8'd33}: color_data = 12'hd21;
			{8'd194, 8'd34}: color_data = 12'hd31;
			{8'd194, 8'd35}: color_data = 12'hd31;
			{8'd194, 8'd36}: color_data = 12'he41;
			{8'd194, 8'd37}: color_data = 12'he41;
			{8'd194, 8'd38}: color_data = 12'hd41;
			{8'd194, 8'd39}: color_data = 12'hd40;
			{8'd194, 8'd47}: color_data = 12'hc70;
			{8'd194, 8'd48}: color_data = 12'hc70;
			{8'd194, 8'd49}: color_data = 12'hc80;
			{8'd194, 8'd50}: color_data = 12'hc80;
			{8'd194, 8'd51}: color_data = 12'hc80;
			{8'd194, 8'd52}: color_data = 12'hb70;
			{8'd194, 8'd53}: color_data = 12'ha60;
			{8'd195, 8'd31}: color_data = 12'hc21;
			{8'd195, 8'd32}: color_data = 12'hd21;
			{8'd195, 8'd33}: color_data = 12'he21;
			{8'd195, 8'd34}: color_data = 12'he31;
			{8'd195, 8'd35}: color_data = 12'he31;
			{8'd195, 8'd36}: color_data = 12'he41;
			{8'd195, 8'd37}: color_data = 12'he41;
			{8'd195, 8'd38}: color_data = 12'hd41;
			{8'd195, 8'd39}: color_data = 12'hc40;
			{8'd195, 8'd47}: color_data = 12'hb71;
			{8'd195, 8'd48}: color_data = 12'ha60;
			{8'd195, 8'd49}: color_data = 12'ha70;
			{8'd195, 8'd50}: color_data = 12'ha70;
			{8'd195, 8'd51}: color_data = 12'h960;
			{8'd195, 8'd52}: color_data = 12'h860;
			{8'd195, 8'd53}: color_data = 12'h770;
			{8'd196, 8'd31}: color_data = 12'hc30;
			{8'd196, 8'd32}: color_data = 12'hd21;
			{8'd196, 8'd33}: color_data = 12'hd21;
			{8'd196, 8'd34}: color_data = 12'hd31;
			{8'd196, 8'd35}: color_data = 12'hd31;
			{8'd196, 8'd36}: color_data = 12'he41;
			{8'd196, 8'd37}: color_data = 12'he41;
			{8'd196, 8'd38}: color_data = 12'hd41;
			{8'd196, 8'd39}: color_data = 12'hf70;
			{8'd203, 8'd33}: color_data = 12'hd02;
			{8'd203, 8'd34}: color_data = 12'hb02;
			{8'd203, 8'd35}: color_data = 12'hb21;
			{8'd203, 8'd36}: color_data = 12'hd20;
			{8'd204, 8'd33}: color_data = 12'hc11;
			{8'd204, 8'd34}: color_data = 12'hd11;
			{8'd204, 8'd35}: color_data = 12'hd11;
			{8'd204, 8'd36}: color_data = 12'hc21;
			{8'd204, 8'd37}: color_data = 12'ha20;
			{8'd204, 8'd43}: color_data = 12'hc71;
			{8'd204, 8'd44}: color_data = 12'he61;
			{8'd204, 8'd45}: color_data = 12'he61;
			{8'd204, 8'd46}: color_data = 12'he61;
			{8'd204, 8'd47}: color_data = 12'hb50;
			{8'd204, 8'd48}: color_data = 12'h850;
			{8'd204, 8'd49}: color_data = 12'h850;
			{8'd204, 8'd50}: color_data = 12'h950;
			{8'd204, 8'd51}: color_data = 12'ha60;
			{8'd204, 8'd52}: color_data = 12'hb70;
			{8'd204, 8'd53}: color_data = 12'hb70;
			{8'd205, 8'd32}: color_data = 12'hf00;
			{8'd205, 8'd33}: color_data = 12'hc11;
			{8'd205, 8'd34}: color_data = 12'hd11;
			{8'd205, 8'd35}: color_data = 12'he21;
			{8'd205, 8'd36}: color_data = 12'hd21;
			{8'd205, 8'd37}: color_data = 12'hb21;
			{8'd205, 8'd38}: color_data = 12'hb31;
			{8'd205, 8'd39}: color_data = 12'ha31;
			{8'd205, 8'd40}: color_data = 12'hc31;
			{8'd205, 8'd41}: color_data = 12'hd51;
			{8'd205, 8'd42}: color_data = 12'hc51;
			{8'd205, 8'd43}: color_data = 12'hc61;
			{8'd205, 8'd44}: color_data = 12'hd61;
			{8'd205, 8'd45}: color_data = 12'hd61;
			{8'd205, 8'd46}: color_data = 12'hd61;
			{8'd205, 8'd47}: color_data = 12'hd70;
			{8'd205, 8'd48}: color_data = 12'hc70;
			{8'd205, 8'd49}: color_data = 12'hb70;
			{8'd205, 8'd50}: color_data = 12'hc70;
			{8'd205, 8'd51}: color_data = 12'hd80;
			{8'd205, 8'd52}: color_data = 12'hd80;
			{8'd205, 8'd53}: color_data = 12'hb80;
			{8'd205, 8'd54}: color_data = 12'h000;
			{8'd206, 8'd32}: color_data = 12'hb01;
			{8'd206, 8'd33}: color_data = 12'hc01;
			{8'd206, 8'd34}: color_data = 12'hd11;
			{8'd206, 8'd35}: color_data = 12'hd21;
			{8'd206, 8'd36}: color_data = 12'hd21;
			{8'd206, 8'd37}: color_data = 12'hd31;
			{8'd206, 8'd38}: color_data = 12'hc31;
			{8'd206, 8'd39}: color_data = 12'hc31;
			{8'd206, 8'd40}: color_data = 12'hd41;
			{8'd206, 8'd41}: color_data = 12'he51;
			{8'd206, 8'd42}: color_data = 12'he51;
			{8'd206, 8'd43}: color_data = 12'he61;
			{8'd206, 8'd44}: color_data = 12'he71;
			{8'd206, 8'd45}: color_data = 12'he71;
			{8'd206, 8'd46}: color_data = 12'he71;
			{8'd206, 8'd47}: color_data = 12'he80;
			{8'd206, 8'd48}: color_data = 12'he80;
			{8'd206, 8'd49}: color_data = 12'he80;
			{8'd206, 8'd50}: color_data = 12'he90;
			{8'd206, 8'd51}: color_data = 12'he90;
			{8'd206, 8'd52}: color_data = 12'he90;
			{8'd206, 8'd53}: color_data = 12'hc80;
			{8'd206, 8'd54}: color_data = 12'h0f0;
			{8'd207, 8'd32}: color_data = 12'hb01;
			{8'd207, 8'd33}: color_data = 12'hc01;
			{8'd207, 8'd34}: color_data = 12'hd11;
			{8'd207, 8'd35}: color_data = 12'hd21;
			{8'd207, 8'd36}: color_data = 12'hd21;
			{8'd207, 8'd37}: color_data = 12'hd31;
			{8'd207, 8'd38}: color_data = 12'he41;
			{8'd207, 8'd39}: color_data = 12'he41;
			{8'd207, 8'd40}: color_data = 12'he51;
			{8'd207, 8'd41}: color_data = 12'he51;
			{8'd207, 8'd42}: color_data = 12'he51;
			{8'd207, 8'd43}: color_data = 12'he61;
			{8'd207, 8'd44}: color_data = 12'he61;
			{8'd207, 8'd45}: color_data = 12'he61;
			{8'd207, 8'd46}: color_data = 12'he71;
			{8'd207, 8'd47}: color_data = 12'he80;
			{8'd207, 8'd48}: color_data = 12'he80;
			{8'd207, 8'd49}: color_data = 12'he80;
			{8'd207, 8'd50}: color_data = 12'he90;
			{8'd207, 8'd51}: color_data = 12'he90;
			{8'd207, 8'd52}: color_data = 12'he90;
			{8'd207, 8'd53}: color_data = 12'hc80;
			{8'd207, 8'd54}: color_data = 12'h000;
			{8'd208, 8'd32}: color_data = 12'hb01;
			{8'd208, 8'd33}: color_data = 12'hc01;
			{8'd208, 8'd34}: color_data = 12'hd11;
			{8'd208, 8'd35}: color_data = 12'hd21;
			{8'd208, 8'd36}: color_data = 12'he21;
			{8'd208, 8'd37}: color_data = 12'hd31;
			{8'd208, 8'd38}: color_data = 12'he41;
			{8'd208, 8'd39}: color_data = 12'he41;
			{8'd208, 8'd40}: color_data = 12'he51;
			{8'd208, 8'd41}: color_data = 12'he51;
			{8'd208, 8'd42}: color_data = 12'he51;
			{8'd208, 8'd43}: color_data = 12'he61;
			{8'd208, 8'd44}: color_data = 12'he61;
			{8'd208, 8'd45}: color_data = 12'he61;
			{8'd208, 8'd46}: color_data = 12'he71;
			{8'd208, 8'd47}: color_data = 12'he80;
			{8'd208, 8'd48}: color_data = 12'hd80;
			{8'd208, 8'd49}: color_data = 12'hd80;
			{8'd208, 8'd50}: color_data = 12'hd80;
			{8'd208, 8'd51}: color_data = 12'hd80;
			{8'd208, 8'd52}: color_data = 12'hd80;
			{8'd208, 8'd53}: color_data = 12'hb70;
			{8'd208, 8'd54}: color_data = 12'h000;
			{8'd209, 8'd32}: color_data = 12'hb01;
			{8'd209, 8'd33}: color_data = 12'hd01;
			{8'd209, 8'd34}: color_data = 12'hd11;
			{8'd209, 8'd35}: color_data = 12'hc11;
			{8'd209, 8'd36}: color_data = 12'hb21;
			{8'd209, 8'd37}: color_data = 12'hb20;
			{8'd209, 8'd38}: color_data = 12'hb31;
			{8'd209, 8'd39}: color_data = 12'hc31;
			{8'd209, 8'd40}: color_data = 12'hb41;
			{8'd209, 8'd41}: color_data = 12'ha41;
			{8'd209, 8'd42}: color_data = 12'hb41;
			{8'd209, 8'd43}: color_data = 12'hd61;
			{8'd209, 8'd44}: color_data = 12'he61;
			{8'd209, 8'd45}: color_data = 12'he61;
			{8'd209, 8'd46}: color_data = 12'he71;
			{8'd209, 8'd47}: color_data = 12'hd70;
			{8'd209, 8'd48}: color_data = 12'hc70;
			{8'd209, 8'd49}: color_data = 12'hb70;
			{8'd209, 8'd50}: color_data = 12'ha60;
			{8'd209, 8'd51}: color_data = 12'ha60;
			{8'd209, 8'd52}: color_data = 12'ha60;
			{8'd209, 8'd53}: color_data = 12'ha60;
			{8'd210, 8'd31}: color_data = 12'h901;
			{8'd210, 8'd32}: color_data = 12'hb01;
			{8'd210, 8'd33}: color_data = 12'hd01;
			{8'd210, 8'd34}: color_data = 12'hd11;
			{8'd210, 8'd35}: color_data = 12'ha11;
			{8'd210, 8'd36}: color_data = 12'h811;
			{8'd210, 8'd37}: color_data = 12'h910;
			{8'd210, 8'd38}: color_data = 12'h711;
			{8'd210, 8'd42}: color_data = 12'ha40;
			{8'd210, 8'd43}: color_data = 12'hd61;
			{8'd210, 8'd44}: color_data = 12'he61;
			{8'd210, 8'd45}: color_data = 12'he61;
			{8'd210, 8'd46}: color_data = 12'hd61;
			{8'd210, 8'd47}: color_data = 12'hb60;
			{8'd210, 8'd48}: color_data = 12'ha50;
			{8'd210, 8'd50}: color_data = 12'hff0;
			{8'd210, 8'd51}: color_data = 12'h930;
			{8'd210, 8'd52}: color_data = 12'h330;
			{8'd211, 8'd31}: color_data = 12'h901;
			{8'd211, 8'd32}: color_data = 12'hb01;
			{8'd211, 8'd33}: color_data = 12'hd01;
			{8'd211, 8'd34}: color_data = 12'hc11;
			{8'd211, 8'd35}: color_data = 12'ha10;
			{8'd211, 8'd42}: color_data = 12'hc50;
			{8'd211, 8'd43}: color_data = 12'hd61;
			{8'd211, 8'd44}: color_data = 12'he61;
			{8'd211, 8'd45}: color_data = 12'he61;
			{8'd211, 8'd46}: color_data = 12'hc60;
			{8'd211, 8'd47}: color_data = 12'h950;
			{8'd212, 8'd31}: color_data = 12'ha01;
			{8'd212, 8'd32}: color_data = 12'hc01;
			{8'd212, 8'd33}: color_data = 12'hd01;
			{8'd212, 8'd34}: color_data = 12'hc11;
			{8'd212, 8'd35}: color_data = 12'h910;
			{8'd212, 8'd42}: color_data = 12'hc51;
			{8'd212, 8'd43}: color_data = 12'hd61;
			{8'd212, 8'd44}: color_data = 12'he61;
			{8'd212, 8'd45}: color_data = 12'he61;
			{8'd212, 8'd46}: color_data = 12'hd61;
			{8'd212, 8'd47}: color_data = 12'hb60;
			{8'd212, 8'd48}: color_data = 12'ha50;
			{8'd213, 8'd31}: color_data = 12'ha01;
			{8'd213, 8'd32}: color_data = 12'hc01;
			{8'd213, 8'd33}: color_data = 12'hd01;
			{8'd213, 8'd34}: color_data = 12'hb11;
			{8'd213, 8'd35}: color_data = 12'h810;
			{8'd213, 8'd42}: color_data = 12'hc51;
			{8'd213, 8'd43}: color_data = 12'he61;
			{8'd213, 8'd44}: color_data = 12'he61;
			{8'd213, 8'd45}: color_data = 12'he61;
			{8'd213, 8'd46}: color_data = 12'he71;
			{8'd213, 8'd47}: color_data = 12'hd70;
			{8'd213, 8'd48}: color_data = 12'hc70;
			{8'd213, 8'd49}: color_data = 12'ha60;
			{8'd213, 8'd50}: color_data = 12'h950;
			{8'd214, 8'd30}: color_data = 12'h901;
			{8'd214, 8'd31}: color_data = 12'hb01;
			{8'd214, 8'd32}: color_data = 12'hd01;
			{8'd214, 8'd33}: color_data = 12'hd01;
			{8'd214, 8'd34}: color_data = 12'hc11;
			{8'd214, 8'd35}: color_data = 12'ha10;
			{8'd214, 8'd36}: color_data = 12'h810;
			{8'd214, 8'd41}: color_data = 12'hb40;
			{8'd214, 8'd42}: color_data = 12'hc51;
			{8'd214, 8'd43}: color_data = 12'he61;
			{8'd214, 8'd44}: color_data = 12'he61;
			{8'd214, 8'd45}: color_data = 12'he61;
			{8'd214, 8'd46}: color_data = 12'he71;
			{8'd214, 8'd47}: color_data = 12'he80;
			{8'd214, 8'd48}: color_data = 12'he80;
			{8'd214, 8'd49}: color_data = 12'hd80;
			{8'd214, 8'd50}: color_data = 12'hb70;
			{8'd214, 8'd51}: color_data = 12'ha60;
			{8'd214, 8'd52}: color_data = 12'h550;
			{8'd215, 8'd30}: color_data = 12'h901;
			{8'd215, 8'd31}: color_data = 12'hb01;
			{8'd215, 8'd32}: color_data = 12'hd01;
			{8'd215, 8'd33}: color_data = 12'hd01;
			{8'd215, 8'd34}: color_data = 12'hd11;
			{8'd215, 8'd35}: color_data = 12'hd11;
			{8'd215, 8'd36}: color_data = 12'ha10;
			{8'd215, 8'd37}: color_data = 12'h810;
			{8'd215, 8'd40}: color_data = 12'ha40;
			{8'd215, 8'd41}: color_data = 12'hc41;
			{8'd215, 8'd42}: color_data = 12'hd51;
			{8'd215, 8'd43}: color_data = 12'he61;
			{8'd215, 8'd44}: color_data = 12'hd61;
			{8'd215, 8'd45}: color_data = 12'hc51;
			{8'd215, 8'd46}: color_data = 12'hb60;
			{8'd215, 8'd47}: color_data = 12'hd70;
			{8'd215, 8'd48}: color_data = 12'he80;
			{8'd215, 8'd49}: color_data = 12'he80;
			{8'd215, 8'd50}: color_data = 12'he90;
			{8'd215, 8'd51}: color_data = 12'hc80;
			{8'd215, 8'd52}: color_data = 12'hb70;
			{8'd215, 8'd53}: color_data = 12'ha60;
			{8'd216, 8'd30}: color_data = 12'h901;
			{8'd216, 8'd31}: color_data = 12'hc02;
			{8'd216, 8'd32}: color_data = 12'hd01;
			{8'd216, 8'd33}: color_data = 12'hd01;
			{8'd216, 8'd34}: color_data = 12'hd11;
			{8'd216, 8'd35}: color_data = 12'hd21;
			{8'd216, 8'd36}: color_data = 12'hc21;
			{8'd216, 8'd37}: color_data = 12'ha21;
			{8'd216, 8'd38}: color_data = 12'h921;
			{8'd216, 8'd39}: color_data = 12'ha21;
			{8'd216, 8'd40}: color_data = 12'hc41;
			{8'd216, 8'd41}: color_data = 12'he51;
			{8'd216, 8'd42}: color_data = 12'he51;
			{8'd216, 8'd43}: color_data = 12'he61;
			{8'd216, 8'd44}: color_data = 12'hc51;
			{8'd216, 8'd45}: color_data = 12'ha41;
			{8'd216, 8'd46}: color_data = 12'h940;
			{8'd216, 8'd47}: color_data = 12'hc60;
			{8'd216, 8'd48}: color_data = 12'he80;
			{8'd216, 8'd49}: color_data = 12'he80;
			{8'd216, 8'd50}: color_data = 12'he90;
			{8'd216, 8'd51}: color_data = 12'he90;
			{8'd216, 8'd52}: color_data = 12'hd80;
			{8'd216, 8'd53}: color_data = 12'hc70;
			{8'd216, 8'd54}: color_data = 12'h960;
			{8'd217, 8'd30}: color_data = 12'h801;
			{8'd217, 8'd31}: color_data = 12'ha01;
			{8'd217, 8'd32}: color_data = 12'hd01;
			{8'd217, 8'd33}: color_data = 12'hd01;
			{8'd217, 8'd34}: color_data = 12'hd11;
			{8'd217, 8'd35}: color_data = 12'hd21;
			{8'd217, 8'd36}: color_data = 12'hd21;
			{8'd217, 8'd37}: color_data = 12'hd31;
			{8'd217, 8'd38}: color_data = 12'hb31;
			{8'd217, 8'd39}: color_data = 12'hc31;
			{8'd217, 8'd40}: color_data = 12'he51;
			{8'd217, 8'd41}: color_data = 12'he51;
			{8'd217, 8'd42}: color_data = 12'hd51;
			{8'd217, 8'd43}: color_data = 12'hb51;
			{8'd217, 8'd44}: color_data = 12'ha41;
			{8'd217, 8'd47}: color_data = 12'hb60;
			{8'd217, 8'd48}: color_data = 12'hd70;
			{8'd217, 8'd49}: color_data = 12'he80;
			{8'd217, 8'd50}: color_data = 12'he90;
			{8'd217, 8'd51}: color_data = 12'he90;
			{8'd217, 8'd52}: color_data = 12'he90;
			{8'd217, 8'd53}: color_data = 12'hc80;
			{8'd217, 8'd54}: color_data = 12'ha70;
			{8'd218, 8'd31}: color_data = 12'h801;
			{8'd218, 8'd32}: color_data = 12'ha01;
			{8'd218, 8'd33}: color_data = 12'hc01;
			{8'd218, 8'd34}: color_data = 12'hd11;
			{8'd218, 8'd35}: color_data = 12'hd21;
			{8'd218, 8'd36}: color_data = 12'hd21;
			{8'd218, 8'd37}: color_data = 12'hd31;
			{8'd218, 8'd38}: color_data = 12'hd31;
			{8'd218, 8'd39}: color_data = 12'he41;
			{8'd218, 8'd40}: color_data = 12'he51;
			{8'd218, 8'd41}: color_data = 12'hd51;
			{8'd218, 8'd42}: color_data = 12'hb41;
			{8'd218, 8'd43}: color_data = 12'h930;
			{8'd218, 8'd47}: color_data = 12'h950;
			{8'd218, 8'd48}: color_data = 12'hb60;
			{8'd218, 8'd49}: color_data = 12'he80;
			{8'd218, 8'd50}: color_data = 12'he90;
			{8'd218, 8'd51}: color_data = 12'he90;
			{8'd218, 8'd52}: color_data = 12'he90;
			{8'd218, 8'd53}: color_data = 12'hd80;
			{8'd218, 8'd54}: color_data = 12'hc80;
			{8'd219, 8'd32}: color_data = 12'h801;
			{8'd219, 8'd33}: color_data = 12'ha01;
			{8'd219, 8'd34}: color_data = 12'hc11;
			{8'd219, 8'd35}: color_data = 12'hd21;
			{8'd219, 8'd36}: color_data = 12'hd21;
			{8'd219, 8'd37}: color_data = 12'hd31;
			{8'd219, 8'd38}: color_data = 12'hd31;
			{8'd219, 8'd39}: color_data = 12'he41;
			{8'd219, 8'd40}: color_data = 12'hd41;
			{8'd219, 8'd41}: color_data = 12'hb40;
			{8'd219, 8'd42}: color_data = 12'h930;
			{8'd219, 8'd47}: color_data = 12'h930;
			{8'd219, 8'd48}: color_data = 12'ha60;
			{8'd219, 8'd49}: color_data = 12'hd80;
			{8'd219, 8'd50}: color_data = 12'he90;
			{8'd219, 8'd51}: color_data = 12'he90;
			{8'd219, 8'd52}: color_data = 12'he90;
			{8'd219, 8'd53}: color_data = 12'hd80;
			{8'd219, 8'd54}: color_data = 12'hc80;
			{8'd220, 8'd33}: color_data = 12'h901;
			{8'd220, 8'd34}: color_data = 12'ha11;
			{8'd220, 8'd35}: color_data = 12'hc11;
			{8'd220, 8'd36}: color_data = 12'hd21;
			{8'd220, 8'd37}: color_data = 12'hd31;
			{8'd220, 8'd38}: color_data = 12'he31;
			{8'd220, 8'd39}: color_data = 12'hd31;
			{8'd220, 8'd40}: color_data = 12'ha30;
			{8'd220, 8'd41}: color_data = 12'h820;
			{8'd220, 8'd48}: color_data = 12'ha60;
			{8'd220, 8'd49}: color_data = 12'hc70;
			{8'd220, 8'd50}: color_data = 12'he90;
			{8'd220, 8'd51}: color_data = 12'he90;
			{8'd220, 8'd52}: color_data = 12'he90;
			{8'd220, 8'd53}: color_data = 12'hd80;
			{8'd220, 8'd54}: color_data = 12'hb70;
			{8'd221, 8'd34}: color_data = 12'h710;
			{8'd221, 8'd35}: color_data = 12'ha11;
			{8'd221, 8'd36}: color_data = 12'hc21;
			{8'd221, 8'd37}: color_data = 12'he31;
			{8'd221, 8'd38}: color_data = 12'hd31;
			{8'd221, 8'd39}: color_data = 12'hb31;
			{8'd221, 8'd40}: color_data = 12'h820;
			{8'd221, 8'd48}: color_data = 12'h550;
			{8'd221, 8'd49}: color_data = 12'hb70;
			{8'd221, 8'd50}: color_data = 12'hd80;
			{8'd221, 8'd51}: color_data = 12'he90;
			{8'd221, 8'd52}: color_data = 12'hd90;
			{8'd221, 8'd53}: color_data = 12'hc80;
			{8'd221, 8'd54}: color_data = 12'ha70;
			{8'd222, 8'd35}: color_data = 12'h400;
			{8'd222, 8'd36}: color_data = 12'ha11;
			{8'd222, 8'd37}: color_data = 12'hc31;
			{8'd222, 8'd38}: color_data = 12'hb31;
			{8'd222, 8'd39}: color_data = 12'h820;
			{8'd222, 8'd49}: color_data = 12'ha60;
			{8'd222, 8'd50}: color_data = 12'hc70;
			{8'd222, 8'd51}: color_data = 12'hd80;
			{8'd222, 8'd52}: color_data = 12'hc80;
			{8'd222, 8'd53}: color_data = 12'hc80;
            default: color_data = 12'h3b9;
        endcase
endmodule   
