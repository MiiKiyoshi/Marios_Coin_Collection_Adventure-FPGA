module coin_rom(
        input wire clk,
        input wire [4:0] x,
        input wire [4:0] y,
        output reg [11:0] color_data
);

    (* rom_style = "block" *)

    //signal declaration
    reg [4:0] x_reg;
    reg [4:0] y_reg;

    always @(posedge clk) begin
        x_reg <= x;
        y_reg <= y;
    end

    always @*
        case ({x_reg, y_reg})
    			// right: 5'd21, bottom: 5'd31
			{5'd0, 5'd0}: color_data = 12'h3b9;
			{5'd0, 5'd1}: color_data = 12'h3b9;
			{5'd0, 5'd2}: color_data = 12'h3b9;
			{5'd0, 5'd3}: color_data = 12'h3b9;
			{5'd0, 5'd4}: color_data = 12'h3b9;
			{5'd0, 5'd5}: color_data = 12'h3b9;
			{5'd0, 5'd6}: color_data = 12'he70;
			{5'd0, 5'd7}: color_data = 12'hf92;
			{5'd0, 5'd8}: color_data = 12'hf93;
			{5'd0, 5'd9}: color_data = 12'hf93;
			{5'd0, 5'd10}: color_data = 12'hf93;
			{5'd0, 5'd11}: color_data = 12'hf93;
			{5'd0, 5'd12}: color_data = 12'hf93;
			{5'd0, 5'd13}: color_data = 12'hf93;
			{5'd0, 5'd14}: color_data = 12'hf93;
			{5'd0, 5'd15}: color_data = 12'hf93;
			{5'd0, 5'd16}: color_data = 12'hf93;
			{5'd0, 5'd17}: color_data = 12'hf93;
			{5'd0, 5'd18}: color_data = 12'hf93;
			{5'd0, 5'd19}: color_data = 12'hf93;
			{5'd0, 5'd20}: color_data = 12'hf93;
			{5'd0, 5'd21}: color_data = 12'hf93;
			{5'd0, 5'd22}: color_data = 12'hf93;
			{5'd0, 5'd23}: color_data = 12'hf93;
			{5'd0, 5'd24}: color_data = 12'hf92;
			{5'd0, 5'd25}: color_data = 12'hf81;
			{5'd0, 5'd26}: color_data = 12'h3b9;
			{5'd0, 5'd27}: color_data = 12'h3b9;
			{5'd0, 5'd28}: color_data = 12'h3b9;
			{5'd0, 5'd29}: color_data = 12'h3b9;
			{5'd0, 5'd30}: color_data = 12'h3b9;
			{5'd0, 5'd31}: color_data = 12'h3b9;
			{5'd1, 5'd0}: color_data = 12'h3b9;
			{5'd1, 5'd1}: color_data = 12'h3b9;
			{5'd1, 5'd2}: color_data = 12'h3b9;
			{5'd1, 5'd3}: color_data = 12'h3b9;
			{5'd1, 5'd4}: color_data = 12'h3b9;
			{5'd1, 5'd5}: color_data = 12'h3b9;
			{5'd1, 5'd6}: color_data = 12'he80;
			{5'd1, 5'd7}: color_data = 12'hf93;
			{5'd1, 5'd8}: color_data = 12'hf93;
			{5'd1, 5'd9}: color_data = 12'hf93;
			{5'd1, 5'd10}: color_data = 12'hf93;
			{5'd1, 5'd11}: color_data = 12'hf93;
			{5'd1, 5'd12}: color_data = 12'hf93;
			{5'd1, 5'd13}: color_data = 12'hf93;
			{5'd1, 5'd14}: color_data = 12'hf93;
			{5'd1, 5'd15}: color_data = 12'hf93;
			{5'd1, 5'd16}: color_data = 12'hf93;
			{5'd1, 5'd17}: color_data = 12'hf93;
			{5'd1, 5'd18}: color_data = 12'hf93;
			{5'd1, 5'd19}: color_data = 12'hf93;
			{5'd1, 5'd20}: color_data = 12'hf93;
			{5'd1, 5'd21}: color_data = 12'hf93;
			{5'd1, 5'd22}: color_data = 12'hf93;
			{5'd1, 5'd23}: color_data = 12'hf93;
			{5'd1, 5'd24}: color_data = 12'hf93;
			{5'd1, 5'd25}: color_data = 12'hf92;
			{5'd1, 5'd26}: color_data = 12'h3b9;
			{5'd1, 5'd27}: color_data = 12'h3b9;
			{5'd1, 5'd28}: color_data = 12'h3b9;
			{5'd1, 5'd29}: color_data = 12'h3b9;
			{5'd1, 5'd30}: color_data = 12'h3b9;
			{5'd1, 5'd31}: color_data = 12'h3b9;
			{5'd2, 5'd0}: color_data = 12'h3b9;
			{5'd2, 5'd1}: color_data = 12'h3b9;
			{5'd2, 5'd2}: color_data = 12'hf92;
			{5'd2, 5'd3}: color_data = 12'hf92;
			{5'd2, 5'd4}: color_data = 12'hf92;
			{5'd2, 5'd5}: color_data = 12'hf92;
			{5'd2, 5'd6}: color_data = 12'hf92;
			{5'd2, 5'd7}: color_data = 12'hf93;
			{5'd2, 5'd8}: color_data = 12'hf93;
			{5'd2, 5'd9}: color_data = 12'hf93;
			{5'd2, 5'd10}: color_data = 12'hf93;
			{5'd2, 5'd11}: color_data = 12'hf93;
			{5'd2, 5'd12}: color_data = 12'hf93;
			{5'd2, 5'd13}: color_data = 12'hf93;
			{5'd2, 5'd14}: color_data = 12'hf93;
			{5'd2, 5'd15}: color_data = 12'hf93;
			{5'd2, 5'd16}: color_data = 12'hf93;
			{5'd2, 5'd17}: color_data = 12'hf93;
			{5'd2, 5'd18}: color_data = 12'hf93;
			{5'd2, 5'd19}: color_data = 12'hf93;
			{5'd2, 5'd20}: color_data = 12'hf93;
			{5'd2, 5'd21}: color_data = 12'hf93;
			{5'd2, 5'd22}: color_data = 12'hf93;
			{5'd2, 5'd23}: color_data = 12'hf93;
			{5'd2, 5'd24}: color_data = 12'hf93;
			{5'd2, 5'd25}: color_data = 12'hf93;
			{5'd2, 5'd26}: color_data = 12'hf92;
			{5'd2, 5'd27}: color_data = 12'hf93;
			{5'd2, 5'd28}: color_data = 12'hf92;
			{5'd2, 5'd29}: color_data = 12'hf92;
			{5'd2, 5'd30}: color_data = 12'h3b9;
			{5'd2, 5'd31}: color_data = 12'h3b9;
			{5'd3, 5'd0}: color_data = 12'h3b9;
			{5'd3, 5'd1}: color_data = 12'h3b9;
			{5'd3, 5'd2}: color_data = 12'hf92;
			{5'd3, 5'd3}: color_data = 12'hfa3;
			{5'd3, 5'd4}: color_data = 12'hf93;
			{5'd3, 5'd5}: color_data = 12'hf93;
			{5'd3, 5'd6}: color_data = 12'hf93;
			{5'd3, 5'd7}: color_data = 12'hf93;
			{5'd3, 5'd8}: color_data = 12'hf93;
			{5'd3, 5'd9}: color_data = 12'hf93;
			{5'd3, 5'd10}: color_data = 12'hf93;
			{5'd3, 5'd11}: color_data = 12'hf93;
			{5'd3, 5'd12}: color_data = 12'hf93;
			{5'd3, 5'd13}: color_data = 12'hf93;
			{5'd3, 5'd14}: color_data = 12'hf93;
			{5'd3, 5'd15}: color_data = 12'hf93;
			{5'd3, 5'd16}: color_data = 12'hf93;
			{5'd3, 5'd17}: color_data = 12'hf93;
			{5'd3, 5'd18}: color_data = 12'hf93;
			{5'd3, 5'd19}: color_data = 12'hf93;
			{5'd3, 5'd20}: color_data = 12'hf93;
			{5'd3, 5'd21}: color_data = 12'hf93;
			{5'd3, 5'd22}: color_data = 12'hf93;
			{5'd3, 5'd23}: color_data = 12'hf93;
			{5'd3, 5'd24}: color_data = 12'hf93;
			{5'd3, 5'd25}: color_data = 12'hf93;
			{5'd3, 5'd26}: color_data = 12'hf93;
			{5'd3, 5'd27}: color_data = 12'hf93;
			{5'd3, 5'd28}: color_data = 12'hfa3;
			{5'd3, 5'd29}: color_data = 12'hf92;
			{5'd3, 5'd30}: color_data = 12'h3b9;
			{5'd3, 5'd31}: color_data = 12'h3b9;
			{5'd4, 5'd0}: color_data = 12'hf82;
			{5'd4, 5'd1}: color_data = 12'hf92;
			{5'd4, 5'd2}: color_data = 12'hf92;
			{5'd4, 5'd3}: color_data = 12'hf93;
			{5'd4, 5'd4}: color_data = 12'hf93;
			{5'd4, 5'd5}: color_data = 12'hf93;
			{5'd4, 5'd6}: color_data = 12'hf93;
			{5'd4, 5'd7}: color_data = 12'hd61;
			{5'd4, 5'd8}: color_data = 12'hd61;
			{5'd4, 5'd9}: color_data = 12'hd61;
			{5'd4, 5'd10}: color_data = 12'hd61;
			{5'd4, 5'd11}: color_data = 12'hd61;
			{5'd4, 5'd12}: color_data = 12'hd61;
			{5'd4, 5'd13}: color_data = 12'hd61;
			{5'd4, 5'd14}: color_data = 12'hd61;
			{5'd4, 5'd15}: color_data = 12'hd61;
			{5'd4, 5'd16}: color_data = 12'hd61;
			{5'd4, 5'd17}: color_data = 12'hd61;
			{5'd4, 5'd18}: color_data = 12'hd61;
			{5'd4, 5'd19}: color_data = 12'hd61;
			{5'd4, 5'd20}: color_data = 12'hd61;
			{5'd4, 5'd21}: color_data = 12'hd61;
			{5'd4, 5'd22}: color_data = 12'hd61;
			{5'd4, 5'd23}: color_data = 12'hd61;
			{5'd4, 5'd24}: color_data = 12'hd61;
			{5'd4, 5'd25}: color_data = 12'hf83;
			{5'd4, 5'd26}: color_data = 12'hf93;
			{5'd4, 5'd27}: color_data = 12'hf93;
			{5'd4, 5'd28}: color_data = 12'hf93;
			{5'd4, 5'd29}: color_data = 12'hf93;
			{5'd4, 5'd30}: color_data = 12'hf92;
			{5'd4, 5'd31}: color_data = 12'hf82;
			{5'd5, 5'd0}: color_data = 12'hf93;
			{5'd5, 5'd1}: color_data = 12'hf93;
			{5'd5, 5'd2}: color_data = 12'hf93;
			{5'd5, 5'd3}: color_data = 12'hf93;
			{5'd5, 5'd4}: color_data = 12'hf93;
			{5'd5, 5'd5}: color_data = 12'hf93;
			{5'd5, 5'd6}: color_data = 12'hf93;
			{5'd5, 5'd7}: color_data = 12'hc40;
			{5'd5, 5'd8}: color_data = 12'hc40;
			{5'd5, 5'd9}: color_data = 12'hc40;
			{5'd5, 5'd10}: color_data = 12'hc40;
			{5'd5, 5'd11}: color_data = 12'hc40;
			{5'd5, 5'd12}: color_data = 12'hc40;
			{5'd5, 5'd13}: color_data = 12'hc40;
			{5'd5, 5'd14}: color_data = 12'hc40;
			{5'd5, 5'd15}: color_data = 12'hc40;
			{5'd5, 5'd16}: color_data = 12'hc40;
			{5'd5, 5'd17}: color_data = 12'hc40;
			{5'd5, 5'd18}: color_data = 12'hc40;
			{5'd5, 5'd19}: color_data = 12'hc40;
			{5'd5, 5'd20}: color_data = 12'hc40;
			{5'd5, 5'd21}: color_data = 12'hc40;
			{5'd5, 5'd22}: color_data = 12'hc40;
			{5'd5, 5'd23}: color_data = 12'hc40;
			{5'd5, 5'd24}: color_data = 12'hc40;
			{5'd5, 5'd25}: color_data = 12'hf82;
			{5'd5, 5'd26}: color_data = 12'hf93;
			{5'd5, 5'd27}: color_data = 12'hf93;
			{5'd5, 5'd28}: color_data = 12'hf93;
			{5'd5, 5'd29}: color_data = 12'hf93;
			{5'd5, 5'd30}: color_data = 12'hf93;
			{5'd5, 5'd31}: color_data = 12'hf93;
			{5'd6, 5'd0}: color_data = 12'hf93;
			{5'd6, 5'd1}: color_data = 12'hf93;
			{5'd6, 5'd2}: color_data = 12'hf93;
			{5'd6, 5'd3}: color_data = 12'hf93;
			{5'd6, 5'd4}: color_data = 12'hf83;
			{5'd6, 5'd5}: color_data = 12'he72;
			{5'd6, 5'd6}: color_data = 12'he72;
			{5'd6, 5'd7}: color_data = 12'hd61;
			{5'd6, 5'd8}: color_data = 12'hd61;
			{5'd6, 5'd9}: color_data = 12'hd61;
			{5'd6, 5'd10}: color_data = 12'hd61;
			{5'd6, 5'd11}: color_data = 12'hd61;
			{5'd6, 5'd12}: color_data = 12'hd61;
			{5'd6, 5'd13}: color_data = 12'hd61;
			{5'd6, 5'd14}: color_data = 12'hd61;
			{5'd6, 5'd15}: color_data = 12'hd61;
			{5'd6, 5'd16}: color_data = 12'hd61;
			{5'd6, 5'd17}: color_data = 12'hd61;
			{5'd6, 5'd18}: color_data = 12'hd61;
			{5'd6, 5'd19}: color_data = 12'hd61;
			{5'd6, 5'd20}: color_data = 12'hd61;
			{5'd6, 5'd21}: color_data = 12'hd61;
			{5'd6, 5'd22}: color_data = 12'hd61;
			{5'd6, 5'd23}: color_data = 12'hd61;
			{5'd6, 5'd24}: color_data = 12'hd61;
			{5'd6, 5'd25}: color_data = 12'ha62;
			{5'd6, 5'd26}: color_data = 12'h952;
			{5'd6, 5'd27}: color_data = 12'hc72;
			{5'd6, 5'd28}: color_data = 12'hf93;
			{5'd6, 5'd29}: color_data = 12'hf93;
			{5'd6, 5'd30}: color_data = 12'hf93;
			{5'd6, 5'd31}: color_data = 12'hf93;
			{5'd7, 5'd0}: color_data = 12'hf93;
			{5'd7, 5'd1}: color_data = 12'hf93;
			{5'd7, 5'd2}: color_data = 12'hf93;
			{5'd7, 5'd3}: color_data = 12'hf93;
			{5'd7, 5'd4}: color_data = 12'he72;
			{5'd7, 5'd5}: color_data = 12'hc40;
			{5'd7, 5'd6}: color_data = 12'hc40;
			{5'd7, 5'd7}: color_data = 12'hf93;
			{5'd7, 5'd8}: color_data = 12'hf93;
			{5'd7, 5'd9}: color_data = 12'hf93;
			{5'd7, 5'd10}: color_data = 12'hf93;
			{5'd7, 5'd11}: color_data = 12'hf93;
			{5'd7, 5'd12}: color_data = 12'hf93;
			{5'd7, 5'd13}: color_data = 12'hf93;
			{5'd7, 5'd14}: color_data = 12'hf93;
			{5'd7, 5'd15}: color_data = 12'hf93;
			{5'd7, 5'd16}: color_data = 12'hf93;
			{5'd7, 5'd17}: color_data = 12'hf93;
			{5'd7, 5'd18}: color_data = 12'hf93;
			{5'd7, 5'd19}: color_data = 12'hf93;
			{5'd7, 5'd20}: color_data = 12'hf93;
			{5'd7, 5'd21}: color_data = 12'hf93;
			{5'd7, 5'd22}: color_data = 12'hf93;
			{5'd7, 5'd23}: color_data = 12'hf93;
			{5'd7, 5'd24}: color_data = 12'hf93;
			{5'd7, 5'd25}: color_data = 12'h321;
			{5'd7, 5'd26}: color_data = 12'h000;
			{5'd7, 5'd27}: color_data = 12'h741;
			{5'd7, 5'd28}: color_data = 12'hf93;
			{5'd7, 5'd29}: color_data = 12'hf93;
			{5'd7, 5'd30}: color_data = 12'hf93;
			{5'd7, 5'd31}: color_data = 12'hf93;
			{5'd8, 5'd0}: color_data = 12'hf93;
			{5'd8, 5'd1}: color_data = 12'hf93;
			{5'd8, 5'd2}: color_data = 12'hf93;
			{5'd8, 5'd3}: color_data = 12'hf93;
			{5'd8, 5'd4}: color_data = 12'he72;
			{5'd8, 5'd5}: color_data = 12'hc40;
			{5'd8, 5'd6}: color_data = 12'hc50;
			{5'd8, 5'd7}: color_data = 12'hf93;
			{5'd8, 5'd8}: color_data = 12'hf93;
			{5'd8, 5'd9}: color_data = 12'hf93;
			{5'd8, 5'd10}: color_data = 12'hf93;
			{5'd8, 5'd11}: color_data = 12'hf93;
			{5'd8, 5'd12}: color_data = 12'hf93;
			{5'd8, 5'd13}: color_data = 12'hf93;
			{5'd8, 5'd14}: color_data = 12'hf93;
			{5'd8, 5'd15}: color_data = 12'hf93;
			{5'd8, 5'd16}: color_data = 12'hf93;
			{5'd8, 5'd17}: color_data = 12'hf93;
			{5'd8, 5'd18}: color_data = 12'hf93;
			{5'd8, 5'd19}: color_data = 12'hf93;
			{5'd8, 5'd20}: color_data = 12'hf93;
			{5'd8, 5'd21}: color_data = 12'hf93;
			{5'd8, 5'd22}: color_data = 12'hf93;
			{5'd8, 5'd23}: color_data = 12'hf93;
			{5'd8, 5'd24}: color_data = 12'hf93;
			{5'd8, 5'd25}: color_data = 12'h321;
			{5'd8, 5'd26}: color_data = 12'h000;
			{5'd8, 5'd27}: color_data = 12'h741;
			{5'd8, 5'd28}: color_data = 12'hf93;
			{5'd8, 5'd29}: color_data = 12'hf93;
			{5'd8, 5'd30}: color_data = 12'hf93;
			{5'd8, 5'd31}: color_data = 12'hf93;
			{5'd9, 5'd0}: color_data = 12'hf93;
			{5'd9, 5'd1}: color_data = 12'hf93;
			{5'd9, 5'd2}: color_data = 12'hf93;
			{5'd9, 5'd3}: color_data = 12'hf93;
			{5'd9, 5'd4}: color_data = 12'he72;
			{5'd9, 5'd5}: color_data = 12'hc40;
			{5'd9, 5'd6}: color_data = 12'hc50;
			{5'd9, 5'd7}: color_data = 12'hf93;
			{5'd9, 5'd8}: color_data = 12'hf93;
			{5'd9, 5'd9}: color_data = 12'hf93;
			{5'd9, 5'd10}: color_data = 12'hf93;
			{5'd9, 5'd11}: color_data = 12'hf93;
			{5'd9, 5'd12}: color_data = 12'hf93;
			{5'd9, 5'd13}: color_data = 12'hf93;
			{5'd9, 5'd14}: color_data = 12'hf93;
			{5'd9, 5'd15}: color_data = 12'hf93;
			{5'd9, 5'd16}: color_data = 12'hf93;
			{5'd9, 5'd17}: color_data = 12'hf93;
			{5'd9, 5'd18}: color_data = 12'hf93;
			{5'd9, 5'd19}: color_data = 12'hf93;
			{5'd9, 5'd20}: color_data = 12'hf93;
			{5'd9, 5'd21}: color_data = 12'hf93;
			{5'd9, 5'd22}: color_data = 12'hf93;
			{5'd9, 5'd23}: color_data = 12'hf93;
			{5'd9, 5'd24}: color_data = 12'hf93;
			{5'd9, 5'd25}: color_data = 12'h321;
			{5'd9, 5'd26}: color_data = 12'h000;
			{5'd9, 5'd27}: color_data = 12'h741;
			{5'd9, 5'd28}: color_data = 12'hf93;
			{5'd9, 5'd29}: color_data = 12'hf93;
			{5'd9, 5'd30}: color_data = 12'hf93;
			{5'd9, 5'd31}: color_data = 12'hf93;
			{5'd10, 5'd0}: color_data = 12'hf93;
			{5'd10, 5'd1}: color_data = 12'hf93;
			{5'd10, 5'd2}: color_data = 12'hf93;
			{5'd10, 5'd3}: color_data = 12'hf93;
			{5'd10, 5'd4}: color_data = 12'he82;
			{5'd10, 5'd5}: color_data = 12'hc40;
			{5'd10, 5'd6}: color_data = 12'hc51;
			{5'd10, 5'd7}: color_data = 12'he83;
			{5'd10, 5'd8}: color_data = 12'he83;
			{5'd10, 5'd9}: color_data = 12'he83;
			{5'd10, 5'd10}: color_data = 12'he83;
			{5'd10, 5'd11}: color_data = 12'he83;
			{5'd10, 5'd12}: color_data = 12'he83;
			{5'd10, 5'd13}: color_data = 12'he83;
			{5'd10, 5'd14}: color_data = 12'he83;
			{5'd10, 5'd15}: color_data = 12'he83;
			{5'd10, 5'd16}: color_data = 12'he83;
			{5'd10, 5'd17}: color_data = 12'he83;
			{5'd10, 5'd18}: color_data = 12'he83;
			{5'd10, 5'd19}: color_data = 12'he83;
			{5'd10, 5'd20}: color_data = 12'he83;
			{5'd10, 5'd21}: color_data = 12'he83;
			{5'd10, 5'd22}: color_data = 12'he83;
			{5'd10, 5'd23}: color_data = 12'he83;
			{5'd10, 5'd24}: color_data = 12'he83;
			{5'd10, 5'd25}: color_data = 12'h421;
			{5'd10, 5'd26}: color_data = 12'h000;
			{5'd10, 5'd27}: color_data = 12'h852;
			{5'd10, 5'd28}: color_data = 12'hf93;
			{5'd10, 5'd29}: color_data = 12'hf93;
			{5'd10, 5'd30}: color_data = 12'hf93;
			{5'd10, 5'd31}: color_data = 12'hf93;
			{5'd11, 5'd0}: color_data = 12'hf92;
			{5'd11, 5'd1}: color_data = 12'hf93;
			{5'd11, 5'd2}: color_data = 12'hf93;
			{5'd11, 5'd3}: color_data = 12'hf93;
			{5'd11, 5'd4}: color_data = 12'hf93;
			{5'd11, 5'd5}: color_data = 12'hf93;
			{5'd11, 5'd6}: color_data = 12'he83;
			{5'd11, 5'd7}: color_data = 12'h210;
			{5'd11, 5'd8}: color_data = 12'h000;
			{5'd11, 5'd9}: color_data = 12'h100;
			{5'd11, 5'd10}: color_data = 12'h100;
			{5'd11, 5'd11}: color_data = 12'h100;
			{5'd11, 5'd12}: color_data = 12'h100;
			{5'd11, 5'd13}: color_data = 12'h100;
			{5'd11, 5'd14}: color_data = 12'h100;
			{5'd11, 5'd15}: color_data = 12'h100;
			{5'd11, 5'd16}: color_data = 12'h100;
			{5'd11, 5'd17}: color_data = 12'h100;
			{5'd11, 5'd18}: color_data = 12'h100;
			{5'd11, 5'd19}: color_data = 12'h100;
			{5'd11, 5'd20}: color_data = 12'h100;
			{5'd11, 5'd21}: color_data = 12'h100;
			{5'd11, 5'd22}: color_data = 12'h100;
			{5'd11, 5'd23}: color_data = 12'h100;
			{5'd11, 5'd24}: color_data = 12'h100;
			{5'd11, 5'd25}: color_data = 12'hb72;
			{5'd11, 5'd26}: color_data = 12'hf93;
			{5'd11, 5'd27}: color_data = 12'hf93;
			{5'd11, 5'd28}: color_data = 12'hf93;
			{5'd11, 5'd29}: color_data = 12'hf93;
			{5'd11, 5'd30}: color_data = 12'hf93;
			{5'd11, 5'd31}: color_data = 12'hf93;
			{5'd12, 5'd0}: color_data = 12'hf93;
			{5'd12, 5'd1}: color_data = 12'hf93;
			{5'd12, 5'd2}: color_data = 12'hf93;
			{5'd12, 5'd3}: color_data = 12'hf93;
			{5'd12, 5'd4}: color_data = 12'hf93;
			{5'd12, 5'd5}: color_data = 12'hf93;
			{5'd12, 5'd6}: color_data = 12'he83;
			{5'd12, 5'd7}: color_data = 12'h100;
			{5'd12, 5'd8}: color_data = 12'h000;
			{5'd12, 5'd9}: color_data = 12'h000;
			{5'd12, 5'd10}: color_data = 12'h000;
			{5'd12, 5'd11}: color_data = 12'h000;
			{5'd12, 5'd12}: color_data = 12'h000;
			{5'd12, 5'd13}: color_data = 12'h000;
			{5'd12, 5'd14}: color_data = 12'h000;
			{5'd12, 5'd15}: color_data = 12'h000;
			{5'd12, 5'd16}: color_data = 12'h000;
			{5'd12, 5'd17}: color_data = 12'h000;
			{5'd12, 5'd18}: color_data = 12'h000;
			{5'd12, 5'd19}: color_data = 12'h000;
			{5'd12, 5'd20}: color_data = 12'h000;
			{5'd12, 5'd21}: color_data = 12'h000;
			{5'd12, 5'd22}: color_data = 12'h000;
			{5'd12, 5'd23}: color_data = 12'h000;
			{5'd12, 5'd24}: color_data = 12'h000;
			{5'd12, 5'd25}: color_data = 12'hc72;
			{5'd12, 5'd26}: color_data = 12'hf93;
			{5'd12, 5'd27}: color_data = 12'hf93;
			{5'd12, 5'd28}: color_data = 12'hf93;
			{5'd12, 5'd29}: color_data = 12'hf93;
			{5'd12, 5'd30}: color_data = 12'hf93;
			{5'd12, 5'd31}: color_data = 12'hf93;
			{5'd13, 5'd0}: color_data = 12'h210;
			{5'd13, 5'd1}: color_data = 12'h210;
			{5'd13, 5'd2}: color_data = 12'ha62;
			{5'd13, 5'd3}: color_data = 12'hf93;
			{5'd13, 5'd4}: color_data = 12'hf93;
			{5'd13, 5'd5}: color_data = 12'hf93;
			{5'd13, 5'd6}: color_data = 12'hf93;
			{5'd13, 5'd7}: color_data = 12'hd72;
			{5'd13, 5'd8}: color_data = 12'hc72;
			{5'd13, 5'd9}: color_data = 12'hd72;
			{5'd13, 5'd10}: color_data = 12'hd72;
			{5'd13, 5'd11}: color_data = 12'hd72;
			{5'd13, 5'd12}: color_data = 12'hd72;
			{5'd13, 5'd13}: color_data = 12'hd72;
			{5'd13, 5'd14}: color_data = 12'hd72;
			{5'd13, 5'd15}: color_data = 12'hd72;
			{5'd13, 5'd16}: color_data = 12'hd72;
			{5'd13, 5'd17}: color_data = 12'hd72;
			{5'd13, 5'd18}: color_data = 12'hd72;
			{5'd13, 5'd19}: color_data = 12'hd72;
			{5'd13, 5'd20}: color_data = 12'hd72;
			{5'd13, 5'd21}: color_data = 12'hd72;
			{5'd13, 5'd22}: color_data = 12'hd72;
			{5'd13, 5'd23}: color_data = 12'hd72;
			{5'd13, 5'd24}: color_data = 12'hd72;
			{5'd13, 5'd25}: color_data = 12'hf93;
			{5'd13, 5'd26}: color_data = 12'hf93;
			{5'd13, 5'd27}: color_data = 12'hf93;
			{5'd13, 5'd28}: color_data = 12'hf93;
			{5'd13, 5'd29}: color_data = 12'hc72;
			{5'd13, 5'd30}: color_data = 12'h210;
			{5'd13, 5'd31}: color_data = 12'h210;
			{5'd14, 5'd0}: color_data = 12'h000;
			{5'd14, 5'd1}: color_data = 12'h000;
			{5'd14, 5'd2}: color_data = 12'h952;
			{5'd14, 5'd3}: color_data = 12'hfa3;
			{5'd14, 5'd4}: color_data = 12'hf93;
			{5'd14, 5'd5}: color_data = 12'hf93;
			{5'd14, 5'd6}: color_data = 12'hf93;
			{5'd14, 5'd7}: color_data = 12'hf93;
			{5'd14, 5'd8}: color_data = 12'hf93;
			{5'd14, 5'd9}: color_data = 12'hf93;
			{5'd14, 5'd10}: color_data = 12'hf93;
			{5'd14, 5'd11}: color_data = 12'hf93;
			{5'd14, 5'd12}: color_data = 12'hf93;
			{5'd14, 5'd13}: color_data = 12'hf93;
			{5'd14, 5'd14}: color_data = 12'hf93;
			{5'd14, 5'd15}: color_data = 12'hf93;
			{5'd14, 5'd16}: color_data = 12'hf93;
			{5'd14, 5'd17}: color_data = 12'hf93;
			{5'd14, 5'd18}: color_data = 12'hf93;
			{5'd14, 5'd19}: color_data = 12'hf93;
			{5'd14, 5'd20}: color_data = 12'hf93;
			{5'd14, 5'd21}: color_data = 12'hf93;
			{5'd14, 5'd22}: color_data = 12'hf93;
			{5'd14, 5'd23}: color_data = 12'hf93;
			{5'd14, 5'd24}: color_data = 12'hf93;
			{5'd14, 5'd25}: color_data = 12'hf93;
			{5'd14, 5'd26}: color_data = 12'hf93;
			{5'd14, 5'd27}: color_data = 12'hf93;
			{5'd14, 5'd28}: color_data = 12'hfa3;
			{5'd14, 5'd29}: color_data = 12'hc72;
			{5'd14, 5'd30}: color_data = 12'h000;
			{5'd14, 5'd31}: color_data = 12'h000;
			{5'd15, 5'd0}: color_data = 12'h000;
			{5'd15, 5'd1}: color_data = 12'h000;
			{5'd15, 5'd2}: color_data = 12'h320;
			{5'd15, 5'd3}: color_data = 12'h531;
			{5'd15, 5'd4}: color_data = 12'h531;
			{5'd15, 5'd5}: color_data = 12'h531;
			{5'd15, 5'd6}: color_data = 12'h631;
			{5'd15, 5'd7}: color_data = 12'hf93;
			{5'd15, 5'd8}: color_data = 12'hf93;
			{5'd15, 5'd9}: color_data = 12'hf93;
			{5'd15, 5'd10}: color_data = 12'hf93;
			{5'd15, 5'd11}: color_data = 12'hf93;
			{5'd15, 5'd12}: color_data = 12'hf93;
			{5'd15, 5'd13}: color_data = 12'hf93;
			{5'd15, 5'd14}: color_data = 12'hf93;
			{5'd15, 5'd15}: color_data = 12'hf93;
			{5'd15, 5'd16}: color_data = 12'hf93;
			{5'd15, 5'd17}: color_data = 12'hf93;
			{5'd15, 5'd18}: color_data = 12'hf93;
			{5'd15, 5'd19}: color_data = 12'hf93;
			{5'd15, 5'd20}: color_data = 12'hf93;
			{5'd15, 5'd21}: color_data = 12'hf93;
			{5'd15, 5'd22}: color_data = 12'hf93;
			{5'd15, 5'd23}: color_data = 12'hf93;
			{5'd15, 5'd24}: color_data = 12'hf93;
			{5'd15, 5'd25}: color_data = 12'h741;
			{5'd15, 5'd26}: color_data = 12'h431;
			{5'd15, 5'd27}: color_data = 12'h531;
			{5'd15, 5'd28}: color_data = 12'h531;
			{5'd15, 5'd29}: color_data = 12'h421;
			{5'd15, 5'd30}: color_data = 12'h000;
			{5'd15, 5'd31}: color_data = 12'h000;
			{5'd16, 5'd0}: color_data = 12'h000;
			{5'd16, 5'd1}: color_data = 12'h000;
			{5'd16, 5'd2}: color_data = 12'h000;
			{5'd16, 5'd3}: color_data = 12'h000;
			{5'd16, 5'd4}: color_data = 12'h000;
			{5'd16, 5'd5}: color_data = 12'h000;
			{5'd16, 5'd6}: color_data = 12'h110;
			{5'd16, 5'd7}: color_data = 12'he93;
			{5'd16, 5'd8}: color_data = 12'hf93;
			{5'd16, 5'd9}: color_data = 12'hf93;
			{5'd16, 5'd10}: color_data = 12'hf93;
			{5'd16, 5'd11}: color_data = 12'hf93;
			{5'd16, 5'd12}: color_data = 12'hf93;
			{5'd16, 5'd13}: color_data = 12'hf93;
			{5'd16, 5'd14}: color_data = 12'hf93;
			{5'd16, 5'd15}: color_data = 12'hf93;
			{5'd16, 5'd16}: color_data = 12'hf93;
			{5'd16, 5'd17}: color_data = 12'hf93;
			{5'd16, 5'd18}: color_data = 12'hf93;
			{5'd16, 5'd19}: color_data = 12'hf93;
			{5'd16, 5'd20}: color_data = 12'hf93;
			{5'd16, 5'd21}: color_data = 12'hf93;
			{5'd16, 5'd22}: color_data = 12'hf93;
			{5'd16, 5'd23}: color_data = 12'hf93;
			{5'd16, 5'd24}: color_data = 12'hf93;
			{5'd16, 5'd25}: color_data = 12'h321;
			{5'd16, 5'd26}: color_data = 12'h000;
			{5'd16, 5'd27}: color_data = 12'h000;
			{5'd16, 5'd28}: color_data = 12'h000;
			{5'd16, 5'd29}: color_data = 12'h000;
			{5'd16, 5'd30}: color_data = 12'h000;
			{5'd16, 5'd31}: color_data = 12'h000;
			{5'd17, 5'd0}: color_data = 12'h000;
			{5'd17, 5'd1}: color_data = 12'h000;
			{5'd17, 5'd2}: color_data = 12'h000;
			{5'd17, 5'd3}: color_data = 12'h000;
			{5'd17, 5'd4}: color_data = 12'h000;
			{5'd17, 5'd5}: color_data = 12'h000;
			{5'd17, 5'd6}: color_data = 12'h100;
			{5'd17, 5'd7}: color_data = 12'h741;
			{5'd17, 5'd8}: color_data = 12'h841;
			{5'd17, 5'd9}: color_data = 12'h841;
			{5'd17, 5'd10}: color_data = 12'h841;
			{5'd17, 5'd11}: color_data = 12'h841;
			{5'd17, 5'd12}: color_data = 12'h841;
			{5'd17, 5'd13}: color_data = 12'h841;
			{5'd17, 5'd14}: color_data = 12'h841;
			{5'd17, 5'd15}: color_data = 12'h841;
			{5'd17, 5'd16}: color_data = 12'h841;
			{5'd17, 5'd17}: color_data = 12'h841;
			{5'd17, 5'd18}: color_data = 12'h841;
			{5'd17, 5'd19}: color_data = 12'h841;
			{5'd17, 5'd20}: color_data = 12'h841;
			{5'd17, 5'd21}: color_data = 12'h841;
			{5'd17, 5'd22}: color_data = 12'h841;
			{5'd17, 5'd23}: color_data = 12'h841;
			{5'd17, 5'd24}: color_data = 12'h841;
			{5'd17, 5'd25}: color_data = 12'h210;
			{5'd17, 5'd26}: color_data = 12'h000;
			{5'd17, 5'd27}: color_data = 12'h000;
			{5'd17, 5'd28}: color_data = 12'h000;
			{5'd17, 5'd29}: color_data = 12'h000;
			{5'd17, 5'd30}: color_data = 12'h000;
			{5'd17, 5'd31}: color_data = 12'h000;
			{5'd18, 5'd0}: color_data = 12'h3b9;
			{5'd18, 5'd1}: color_data = 12'h3b9;
			{5'd18, 5'd2}: color_data = 12'h000;
			{5'd18, 5'd3}: color_data = 12'h000;
			{5'd18, 5'd4}: color_data = 12'h000;
			{5'd18, 5'd5}: color_data = 12'h000;
			{5'd18, 5'd6}: color_data = 12'h000;
			{5'd18, 5'd7}: color_data = 12'h000;
			{5'd18, 5'd8}: color_data = 12'h000;
			{5'd18, 5'd9}: color_data = 12'h000;
			{5'd18, 5'd10}: color_data = 12'h000;
			{5'd18, 5'd11}: color_data = 12'h000;
			{5'd18, 5'd12}: color_data = 12'h000;
			{5'd18, 5'd13}: color_data = 12'h000;
			{5'd18, 5'd14}: color_data = 12'h000;
			{5'd18, 5'd15}: color_data = 12'h000;
			{5'd18, 5'd16}: color_data = 12'h000;
			{5'd18, 5'd17}: color_data = 12'h000;
			{5'd18, 5'd18}: color_data = 12'h000;
			{5'd18, 5'd19}: color_data = 12'h000;
			{5'd18, 5'd20}: color_data = 12'h000;
			{5'd18, 5'd21}: color_data = 12'h000;
			{5'd18, 5'd22}: color_data = 12'h000;
			{5'd18, 5'd23}: color_data = 12'h000;
			{5'd18, 5'd24}: color_data = 12'h000;
			{5'd18, 5'd25}: color_data = 12'h000;
			{5'd18, 5'd26}: color_data = 12'h000;
			{5'd18, 5'd27}: color_data = 12'h000;
			{5'd18, 5'd28}: color_data = 12'h000;
			{5'd18, 5'd29}: color_data = 12'h000;
			{5'd18, 5'd30}: color_data = 12'h3b9;
			{5'd18, 5'd31}: color_data = 12'h3b9;
			{5'd19, 5'd0}: color_data = 12'h3b9;
			{5'd19, 5'd1}: color_data = 12'h3b9;
			{5'd19, 5'd2}: color_data = 12'h000;
			{5'd19, 5'd3}: color_data = 12'h000;
			{5'd19, 5'd4}: color_data = 12'h000;
			{5'd19, 5'd5}: color_data = 12'h000;
			{5'd19, 5'd6}: color_data = 12'h000;
			{5'd19, 5'd7}: color_data = 12'h000;
			{5'd19, 5'd8}: color_data = 12'h000;
			{5'd19, 5'd9}: color_data = 12'h000;
			{5'd19, 5'd10}: color_data = 12'h000;
			{5'd19, 5'd11}: color_data = 12'h000;
			{5'd19, 5'd12}: color_data = 12'h000;
			{5'd19, 5'd13}: color_data = 12'h000;
			{5'd19, 5'd14}: color_data = 12'h000;
			{5'd19, 5'd15}: color_data = 12'h000;
			{5'd19, 5'd16}: color_data = 12'h000;
			{5'd19, 5'd17}: color_data = 12'h000;
			{5'd19, 5'd18}: color_data = 12'h000;
			{5'd19, 5'd19}: color_data = 12'h000;
			{5'd19, 5'd20}: color_data = 12'h000;
			{5'd19, 5'd21}: color_data = 12'h000;
			{5'd19, 5'd22}: color_data = 12'h000;
			{5'd19, 5'd23}: color_data = 12'h000;
			{5'd19, 5'd24}: color_data = 12'h000;
			{5'd19, 5'd25}: color_data = 12'h000;
			{5'd19, 5'd26}: color_data = 12'h000;
			{5'd19, 5'd27}: color_data = 12'h000;
			{5'd19, 5'd28}: color_data = 12'h000;
			{5'd19, 5'd29}: color_data = 12'h000;
			{5'd19, 5'd30}: color_data = 12'h3b9;
			{5'd19, 5'd31}: color_data = 12'h3b9;
			{5'd20, 5'd0}: color_data = 12'h3b9;
			{5'd20, 5'd1}: color_data = 12'h3b9;
			{5'd20, 5'd2}: color_data = 12'h3b9;
			{5'd20, 5'd3}: color_data = 12'h3b9;
			{5'd20, 5'd4}: color_data = 12'h3b9;
			{5'd20, 5'd5}: color_data = 12'h3b9;
			{5'd20, 5'd6}: color_data = 12'h000;
			{5'd20, 5'd7}: color_data = 12'h000;
			{5'd20, 5'd8}: color_data = 12'h000;
			{5'd20, 5'd9}: color_data = 12'h000;
			{5'd20, 5'd10}: color_data = 12'h000;
			{5'd20, 5'd11}: color_data = 12'h000;
			{5'd20, 5'd12}: color_data = 12'h000;
			{5'd20, 5'd13}: color_data = 12'h000;
			{5'd20, 5'd14}: color_data = 12'h000;
			{5'd20, 5'd15}: color_data = 12'h000;
			{5'd20, 5'd16}: color_data = 12'h000;
			{5'd20, 5'd17}: color_data = 12'h000;
			{5'd20, 5'd18}: color_data = 12'h000;
			{5'd20, 5'd19}: color_data = 12'h000;
			{5'd20, 5'd20}: color_data = 12'h000;
			{5'd20, 5'd21}: color_data = 12'h000;
			{5'd20, 5'd22}: color_data = 12'h000;
			{5'd20, 5'd23}: color_data = 12'h000;
			{5'd20, 5'd24}: color_data = 12'h000;
			{5'd20, 5'd25}: color_data = 12'h000;
			{5'd20, 5'd26}: color_data = 12'h3b9;
			{5'd20, 5'd27}: color_data = 12'h3b9;
			{5'd20, 5'd28}: color_data = 12'h3b9;
			{5'd20, 5'd29}: color_data = 12'h3b9;
			{5'd20, 5'd30}: color_data = 12'h3b9;
			{5'd20, 5'd31}: color_data = 12'h3b9;
			{5'd21, 5'd0}: color_data = 12'h3b9;
			{5'd21, 5'd1}: color_data = 12'h3b9;
			{5'd21, 5'd2}: color_data = 12'h3b9;
			{5'd21, 5'd3}: color_data = 12'h3b9;
			{5'd21, 5'd4}: color_data = 12'h3b9;
			{5'd21, 5'd5}: color_data = 12'h3b9;
			{5'd21, 5'd6}: color_data = 12'h000;
			{5'd21, 5'd7}: color_data = 12'h000;
			{5'd21, 5'd8}: color_data = 12'h000;
			{5'd21, 5'd9}: color_data = 12'h000;
			{5'd21, 5'd10}: color_data = 12'h000;
			{5'd21, 5'd11}: color_data = 12'h000;
			{5'd21, 5'd12}: color_data = 12'h000;
			{5'd21, 5'd13}: color_data = 12'h000;
			{5'd21, 5'd14}: color_data = 12'h000;
			{5'd21, 5'd15}: color_data = 12'h000;
			{5'd21, 5'd16}: color_data = 12'h000;
			{5'd21, 5'd17}: color_data = 12'h000;
			{5'd21, 5'd18}: color_data = 12'h000;
			{5'd21, 5'd19}: color_data = 12'h000;
			{5'd21, 5'd20}: color_data = 12'h000;
			{5'd21, 5'd21}: color_data = 12'h000;
			{5'd21, 5'd22}: color_data = 12'h000;
			{5'd21, 5'd23}: color_data = 12'h000;
			{5'd21, 5'd24}: color_data = 12'h000;
			{5'd21, 5'd25}: color_data = 12'h000;
			{5'd21, 5'd26}: color_data = 12'h3b9;
			{5'd21, 5'd27}: color_data = 12'h3b9;
			{5'd21, 5'd28}: color_data = 12'h3b9;
			{5'd21, 5'd29}: color_data = 12'h3b9;
			{5'd21, 5'd30}: color_data = 12'h3b9;
			{5'd21, 5'd31}: color_data = 12'h3b9;
            default: color_data = 12'h3b9;
        endcase
endmodule
